Vim�UnDo� Vo��6!�p���Vqs]?������MV?y�6   F   	endmodule   F   	      A       A   A   A    c��    _�                    "        ����                                                                                                                                                                                                                                                                                                                                                             c�     �   "   '   9    �   "   #   9    5�_�                    "        ����                                                                                                                                                                                                                                                                                                                                                             c�     �   !   #   >           �   "   $   >          �   "   $   =    5�_�                    $   	    ����                                                                                                                                                                                                                                                                                                                                                             c�R     �   #   %   =      	next_row_reg = btn_reg_row++;5�_�                    $       ����                                                                                                                                                                                                                                                                                                                                                             c�Y     �   #   %   =      	next_col_reg = btn_reg_row++;5�_�                    $       ����                                                                                                                                                                                                                                                                                                                                                             c�_     �   #   %   =      	next_col_reg = btn_reg_col++;5�_�                    %        ����                                                                                                                                                                                                                                                                                                                                                             c�o     �   %   .   =    �   %   &   =    5�_�      	              &        ����                                                                                                                                                                                                                                                                                                                                                             c�q     �   %   (   E      	begin5�_�      
           	   &        ����                                                                                                                                                                                                                                                                                                                                                             c�s     �   %   '   F       5�_�   	              
   (       ����                                                                                                                                                                                                                                                                                                                                                             c��     �   '   )   F      	next_row_reg = btn_reg_row++;5�_�   
                 *       ����                                                                                                                                                                                                                                                                                                                                                             c��     �   )   +   F      (if (btn_data == 0x4 && btn_reg_col != 0)5�_�                    *   '    ����                                                                                                                                                                                                                                                                                                                                                             c��     �   )   +   F      (if (btn_data == 0x1 && btn_reg_col != 0)5�_�                    *   %    ����                                                                                                                                                                                                                                                                                                                                                             c��     �   )   +   F      ,if (btn_data == 0x1 && btn_reg_col != 0x1DF)5�_�                    "   %    ����                                                                                                                                                                                                                                                                                                                                                             c��     �   !   #   F      (if (btn_data == 0x4 && btn_reg_col != 0)5�_�                       %    ����                                                                                                                                                                                                                                                                                                                                                             c��     �         F      (if (btn_data == 0x8 && btn_reg_row != 0)5�_�                    &   %    ����                                                                                                                                                                                                                                                                                                                                                             c��     �   %   '   F      ,if (btn_data == 0x2 && btn_reg_col != 0x27F)5�_�                    (       ����                                                                                                                                                                                                                                                                                                                                                             c�     �   '   )   F      	next_row_reg = btn_reg_row--;5�_�                    (       ����                                                                                                                                                                                                                                                                                                                                                             c�     �   '   )   F      	next_row_reg = btn_reg_col--;5�_�                    *   "    ����                                                                                                                                                                                                                                                                                                                                                             c�$     �   )   +   F      +if (btn_data == 0x1 && btn_reg_col < 0x1DF)5�_�                    ,       ����                                                                                                                                                                                                                                                                                                                                                             c�(     �   +   -   F      	next_col_reg = btn_reg_col--;5�_�                    -       ����                                                                                                                                                                                                                                                                                                                                                             c�G     �   ,   /   F      	end5�_�                    7       ����                                                                                                                                                                                                                                                                                                                                                             c�e     �   6   9   G      	else begin5�_�                    8        ����                                                                                                                                                                                                                                                                                                                                                             c퉛     �   7   =   H       5�_�                    8       ����                                                                                                                                                                                                                                                                                                                                                             c퉟     �   7   :   L              5�_�                    7       ����                                                                                                                                                                                                                                                                                                                                                             c��     �   6   9   M      	else begin5�_�                    8       ����                                                                                                                                                                                                                                                                                                                                                             c��     �   6   8   N      	else    begin�   7   9   N      	    begin5�_�                    :        ����                                                                                                                                                                                                                                                                                                                                                             c��     �   9   ;   M       5�_�                    7       ����                                                                                                                                                                                                                                                                                                                                                             c�      �   6   9   M      	else begin5�_�                    ;       ����                                                                                                                                                                                                                                                                                                                                                             c�.     �   :   =   N          end5�_�                    <       ����                                                                                                                                                                                                                                                                                                                                                             c�3     �   <   >   O    �   <   =   O    5�_�                     <       ����                                                                                                                                                                                                                                                                                                                                                             c�8     �   :   <   P          end     �   ;   =   P              5�_�      !               8        ����                                                                                                                                                                                                                                                                                                                                                             c�f     �   8   :   O    �   8   9   O    5�_�       "           !   8        ����                                                                                                                                                                                                                                                                                                                                                             c�h     �   7   8           5�_�   !   #           "   8       ����                                                                                                                                                                                                                                                                                                                                                             c�n     �   7   :   O      	   case (btn_m2s_adr_i[5:2])5�_�   "   $           #   9        ����                                                                                                                                                                                                                                                                                                                                                             c�q     �   7   :   P      	   case (btn_m2s_adr_i[5:2])    �   8   :   P       5�_�   #   %           $   :       ����                                                                                                                                                                                                                                                                                                                                                             c�{     �   8   :   P                 1:   btn_reg_row <= next_row_reg;�   9   ;   P      $        btn_reg_row <= next_row_reg;5�_�   $   &           %   :       ����                                                                                                                                                                                                                                                                                                                                                             c튋     �   9   ;   O      $        btn_reg_col <= next_col_reg;5�_�   %   '           &   <       ����                                                                                                                                                                                                                                                                                                                                                             c튕     �   9   <   N      *           2: btn_reg_col <= next_col_reg;    �   :   <   O      	    end      �   ;   =   O      	   case (btn_m2s_adr_i[5:2])5�_�   &   (           '   A       ����                                                                                                                                                                                                                                                                                                                                                             c튯     �   >   @   M      	   case (btn_m2s_adr_i[5:2])    �   ?   A   N      	   	1: btn_reg_row <=     �   @   B   N      	5�_�   '   )           (   9       ����                                                                                                                                                                                                                                                                                                                                                             c�{     �   8   :   L      *           1: btn_reg_row <= next_row_reg;5�_�   (   *           )   9       ����                                                                                                                                                                                                                                                                                                                                                             c틛     �   9   ;   L    �   9   :   L    5�_�   )   +           *   :       ����                                                                                                                                                                                                                                                                                                                                                             c틟     �   8   :   M      4           1: btn_reg_row <= btn_ack_ffnext_row_reg;   ,  btn_reg = btn_ack_ff ? btn_data : btn_reg;�   9   ;   M      /	    btn_reg = btn_ack_ff ? btn_data : btn_reg;5�_�   *   ,           +   9       ����                                                                                                                                                                                                                                                                                                                                                             c틤     �   8   :   L      I           1: btn_reg_row <=   btn_reg = btn_ack_ff ? btn_data : btn_reg;5�_�   +   -           ,   9   &    ����                                                                                                                                                                                                                                                                                                                                                             c틦     �   8   :   L      G           1: btn_reg_row <= btn_reg = btn_ack_ff ? btn_data : btn_reg;5�_�   ,   .           -   9       ����                                                                                                                                                                                                                                                                                                                                                             c틪     �   8   :   L      >           1: btn_reg_row <=  btn_ack_ff ? btn_data : btn_reg;5�_�   -   /           .   9   2    ����                                                                                                                                                                                                                                                                                                                                                             c틲     �   8   :   L      =           1: btn_reg_row <= btn_ack_ff ? btn_data : btn_reg;5�_�   .   0           /   9   .    ����                                                                                                                                                                                                                                                                                                                                                             c��     �   8   :   L      9           1: btn_reg_row <= btn_ack_ff ? next : btn_reg;5�_�   /   1           0   9   @    ����                                                                                                                                                                                                                                                                                                                                                             c��     �   8   :   L      A           1: btn_reg_row <= btn_ack_ff ? next_row_reg : btn_reg;5�_�   0   2           1   :   *    ����                                                                                                                                                                                                                                                                                                                                                             c��     �   9   ;   L      *           2: btn_reg_col <= next_col_reg;5�_�   1   3           2   :       ����                                                                                                                                                                                                                                                                                                                                                             c��     �   9   ;   L                 2: btn_reg_col <= �   :   ;   L    5�_�   2   4           3   :   2    ����                                                                                                                                                                                                                                                                                                                                                             c��     �   9   ;   L      E           2: btn_reg_col <= btn_ack_ff ? next_row_reg : btn_reg_row;5�_�   3   5           4   :   D    ����                                                                                                                                                                                                                                                                                                                                                             c��     �   9   ;   L      E           2: btn_reg_col <= btn_ack_ff ? next_col_reg : btn_reg_row;5�_�   4   6           5   @        ����                                                                                                                                                                                                                                                                                                                                                             c��     �   ?   @          /	    btn_reg = btn_ack_ff ? btn_data : btn_reg;5�_�   5   7           6   <        ����                                                                                                                                                                                                                                                                                                                                                             c��     �   ;   <           5�_�   6   8           7   <        ����                                                                                                                                                                                                                                                                                                                                                             c��     �   ;   <           5�_�   7   9           8   <        ����                                                                                                                                                                                                                                                                                                                                                             c��     �   ;   <           5�_�   8   :           9   <       ����                                                                                                                                                                                                                                                                                                                                                             c��     �   ;   <          	  5�_�   9   =           :   <        ����                                                                                                                                                                                                                                                                                                                                                             c��     �   ;   <          		5�_�   :   >   <       =   B       ����                                                                                                                                                                                                                                                                                                                                                             c�(     �   A   C   F      assign btn_s2m_dat_o = btn_reg;5�_�   =   ?           >   B   -    ����                                                                                                                                                                                                                                                                                                                                                             c�H     �   A   C   F      6assign btn_s2m_dat_o = (btn_m2s_adr_i[5:2]==1)btn_reg;5�_�   >   @           ?   B   .    ����                                                                                                                                                                                                                                                                                                                                                             c�J     �   A   C   F      6assign btn_s2m_dat_o = (btn_m2s_adr_i[5:2]==1)btn_reg;5�_�   ?   A           @   B   8    ����                                                                                                                                                                                                                                                                                                                                                             c�O     �   A   C   F      9assign btn_s2m_dat_o = (btn_m2s_adr_i[5:2]==1) ? btn_reg;5�_�   @               A   F   	    ����                                                                                                                                                                                                                                                                                                                                                             c��    �   E              	endmodule5�_�   :       ;   =   <   B       ����                                                                                                                                                                                                                                                                                                                                                             c�      �   B   C   F    �   A   C   F       assign btn_s2m_dat_o = b(tn_reg;5�_�   :           <   ;   B       ����                                                                                                                                                                                                                                                                                                                                                             c�     �   B   C   F    �   A   C   F       assign btn_s2m_dat_o = (btn_reg;5�_�                     !       ����                                                                                                                                                                                                                                                                                                                                                             c�
     �   !   "   9    �   !   "   9      	begin   	next_row_reg = btn_reg_row++;   	end    5��