Vim�UnDo� z�A�_S���4���]�eB+�d� x��M  f   !        if (sprite_column > 560)   9                          d��    _�                     9       ����                                                                                                                                                                                                                                                                                                                                                             d��    �  8  :  f      !        if (sprite_column > 560) 5��