Vim�UnDo� ��W����Stf�4�S!�wRt�c��gC-1E�      // implementatio   	        #      #  #  #    d
j    _�                            ����                                                                                                                                                                                                                                                                                                                                                             d
J�     �         =    �         =    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d
J�     �         ?      logic   [11:0]      alien2_row;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d
J�     �         ?      logic   [11:0]      alien2_col;5�_�                    	   
    ����                                                                                                                                                                                                                                                                                                                                                             d
J�     �      
   ?           input wire              clk,5�_�                    
   
    ����                                                                                                                                                                                                                                                                                                                                                             d
K      �   	      ?      "    input wire              rst_i,5�_�                       
    ����                                                                                                                                                                                                                                                                                                                                                             d
K      �   
      ?      #    input wire              enable,5�_�                       
    ����                                                                                                                                                                                                                                                                                                                                                             d
K     �   
      ?          input enable,5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             d
K     �   
             #    input logic             enable,5�_�      
           	   
       ����                                                                                                                                                                                                                                                                                                                                                             d
K     �   	   
              input rst_i,5�_�   	              
   	   
    ����                                                                                                                                                                                                                                                                                                                                                             d
K     �      
   =          input clk,5�_�   
                 	   #    ����                                                                                                                                                                                                                                                                                                                                                             d
K     �      
   =      #    input logic                clk,5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             d
K     �   	      =      #	output wire  [3:0]	    alien2_pix,5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             d
K      �   	      =      #	output wire  [3:0]	    alien2_pix,5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             d
K$     �   	      =      %	output wire    [3:0]	    alien2_pix,5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             d
K)     �   	   
          $	output wire    [3:0]	   alien2_pix,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
K/     �         <    �         <    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d
K4     �         =      $	output wire    [3:0]	   alien2_pix,5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d
K6     �         =      !	output wire    [3:0]	   alien2_,5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                             d
K<     �   
      =      *    output logic   [11:0]      alien2_col;5�_�                    
   *    ����                                                                                                                                                                                                                                                                                                                                                             d
K>     �   	      =      *    output logic   [11:0]      alien2_row;5�_�                       )    ����                                                                                                                                                                                                                                                                                                                                                             d
K@     �   
      =      )    output logic   [11:0]      alien2_col5�_�                       '    ����                                                                                                                                                                                                                                                                                                                                                             d
KH     �         =      '	output wire    [3:0]	   alien2_output,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
KM     �         >      '	output wire    [3:0]	   alien2_output,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
KR     �         >          output 5�_�                    	   
    ����                                                                                                                                                                                                                                                                                                                                                             d
KY     �      
   >      (    input logic                clk, rst,5�_�                    	        ����                                                                                                                                                                                                                                                                                                                                                             d
Ke     �      
   >      )    input  logic                clk, rst,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
Kl     �         >          output logic5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
Ky     �         >      logic   [11:0]      alien2_row;5�_�                       !    ����                                                                                                                                                                                                                                                                                                                                                             d
K}     �         >      "logic   [11:0]      alien2_row_ff;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
K�     �         >      logic   [11:0]      alien2_col;5�_�                        &    ����                                                                                                                                                                                                                                                                                                                                                             d
K�     �         >      &logic   [11:0]      alien2_column_reg;5�_�      !                       ����                                                                                                                                                                                                                                                                                                                                                             d
K�     �                alien2_pix = 0;5�_�       "           !           ����                                                                                                                                                                                                                                                                                                                                                             d
K�     �                counter = 0;5�_�   !   #           "           ����                                                                                                                                                                                                                                                                                                                                                             d
K�     �         =      end5�_�   "   $           #           ����                                                                                                                                                                                                                                                                                                                                                             d
K�     �         >       5�_�   #   %           $           ����                                                                                                                                                                                                                                                                                                                                                             d
L     �                clk_wiz_0  clock_divider(   	.clk_in1    (vga_fast_clk),   	.reset      (rst_core),   	.clk_31_5   (vga_31_5_clk));   */5�_�   $   &           %           ����                                                                                                                                                                                                                                                                                                                                                             d
L     �                /*5�_�   %   '           &           ����                                                                                                                                                                                                                                                                                                                                                             d
L	     �                 5�_�   &   (           '           ����                                                                                                                                                                                                                                                                                                                                                             d
L
    �                 5�_�   '   )           (   &        ����                                                                                                                                                                                                                                                                                                                                                             d
L�     �   %   @   6       5�_�   (   *           )   E        ����                                                                                                                                                                                                                                                                                                                                                             d
L�     �   D   E       
            vga_g_reg <= vga_output;            vga_b_reg <= vga_output;           end       else              begin            vga_r_reg <= 4'b0000;           vga_g_reg <= 4'b0000;           vga_b_reg <= 4'b0000;           end           end        5�_�   )   +           *   @        ����                                                                                                                                                                                                                                                                                                                                                             d
L�     �   ?   @          "always_ff @ (posedge vga_31_5_clk)5�_�   *   ,           +   @        ����                                                                                                                                                                                                                                                                                                                                                             d
L�     �   ?   @          begin5�_�   +   -           ,   @       ����                                                                                                                                                                                                                                                                                                                                                             d
L�     �   ?   @              if (video_on)5�_�   ,   .           -   @       ����                                                                                                                                                                                                                                                                                                                                                             d
L�     �   ?   @                  begin5�_�   -   /           .   @       ����                                                                                                                                                                                                                                                                                                                                                             d
L�     �   ?   @                   vga_r_reg <= vga_output;5�_�   .   0           /   '       ����                                                                                                                                                                                                                                                                                                                                                             d
L�     �   &   (   @      , 61 always_ff @ (posedge clk or posedge rst)5�_�   /   1           0   '       ����                                                                                                                                                                                                                                                                                                                                                             d
L�     �   &   (   @      + 6 always_ff @ (posedge clk or posedge rst)5�_�   0   2           1   '       ����                                                                                                                                                                                                                                                                                                                                                             d
L�     �   &   (   @      * 6always_ff @ (posedge clk or posedge rst)5�_�   1   3           2   (       ����                                                                                                                                                                                                                                                                                                                                                             d
L�     �   '   )   @      	 62 begin5�_�   2   4           3   (       ����                                                                                                                                                                                                                                                                                                                                                             d
L�     �   '   )   @       begin5�_�   3   5           4   )       ����                                                                                                                                                                                                                                                                                                                                                             d
M      �   '   *   @      begin        if (rst)�   (   *   @       63     if (rst)5�_�   4   6           5   *       ����                                                                                                                                                                                                                                                                                                                                                             d
M     �   (   +   @          if (rst)            begin�   )   +   @       64         begin5�_�   5   7           6   +       ����                                                                                                                                                                                                                                                                                                                                                             d
M     �   )   ,   @      	    begin            btn_row_ff <= 0;�   *   ,   @       65         btn_row_ff <= 0;5�_�   6   8           7   ,       ����                                                                                                                                                                                                                                                                                                                                                             d
M     �   *   ,   @              btn_row_ff <= 0;            btn_column_ff <= 0;�   +   -   @       66         btn_column_ff <= 0;5�_�   7   9           8   +       ����                                                                                                                                                                                                                                                                                                                                                             d
M     �   *   -   ?      4        btn_row_ff <= 0;         btn_column_ff <= 0;5�_�   8   :           9   -       ����                                                                                                                                                                                                                                                                                                                                                             d
M     �   ,   .   @       67         sprite_row_ff <= 0;5�_�   9   ;           :   .       ����                                                                                                                                                                                                                                                                                                                                                             d
M     �   -   /   @      " 68         sprite_column_ff <= 0;5�_�   :   <           ;   /       ����                                                                                                                                                                                                                                                                                                                                                             d
M     �   -   0   @              sprite_column_ff <= 0;            player_pix_reg <= 0;�   .   0   @        69         player_pix_reg <= 0;5�_�   ;   =           <   -       ����                                                                                                                                                                                                                                                                                                                                                             d
M     �   ,   .   @               sprite_row_ff <= 0;5�_�   <   >           =   0       ����                                                                                                                                                                                                                                                                                                                                                             d
M     �   .   1   @              player_pix_reg <= 0;   `         end                                                                                    �   /   1   @      c 70         end                                                                                    5�_�   =   ?           >   1       ����                                                                                                                                                                                                                                                                                                                                                             d
M     �   0   2   @       71     else5�_�   >   @           ?   2       ����                                                                                                                                                                                                                                                                                                                                                             d
M"     �   0   3   @          else            begin�   1   3   @       72         begin5�_�   ?   A           @   0       ����                                                                                                                                                                                                                                                                                                                                                             d
M)     �   /   1   @      _        end                                                                                    5�_�   @   B           A   3       ����                                                                                                                                                                                                                                                                                                                                                             d
M0     �   1   4   @      	    begin            btn_row_ff <= btn_row;�   2   4   @      " 73         btn_row_ff <= btn_row;5�_�   A   C           B   4       ����                                                                                                                                                                                                                                                                                                                                                             d
M4     �   3   5   @      ( 74         btn_column_ff <= btn_column;5�_�   B   D           C   5       ����                                                                                                                                                                                                                                                                                                                                                             d
M6     �   4   6   @      ( 75         sprite_row_ff <= btn_row_ff;5�_�   C   E           D   6       ����                                                                                                                                                                                                                                                                                                                                                             d
M7     �   5   7   @      . 76         sprite_column_ff <= btn_column_ff;5�_�   D   F           E   7       ����                                                                                                                                                                                                                                                                                                                                                             d
M9     �   6   8   @      ) 77         player_pix_reg <= player_pix;5�_�   E   G           F   8       ����                                                                                                                                                                                                                                                                                                                                                             d
M:     �   6   9   @      &         player_pix_reg <= player_pix;            end�   7   9   @       78         end5�_�   F   H           G   9       ����                                                                                                                                                                                                                                                                                                                                                             d
M>     �   8   :   @       79 end5�_�   G   I           H   :       ����                                                                                                                                                                                                                                                                                                                                                             d
M@     �   8   :   @       end     �   9   ;   @       80  5�_�   H   J           I   :       ����                                                                                                                                                                                                                                                                                                                                                             d
MB     �   9   ;   ?      * 81 assign player_output = player_pix_reg;5�_�   I   K           J   ;       ����                                                                                                                                                                                                                                                                                                                                                             d
MD     �   :   <   ?      & 82 assign player_row = sprite_row_ff;5�_�   J   L           K   <       ����                                                                                                                                                                                                                                                                                                                                                             d
ME     �   ;   =   ?      , 83 assign player_column = sprite_column_ff;5�_�   K   M           L   =       ����                                                                                                                                                                                                                                                                                                                                                             d
MG     �   <   >   ?      " 84 assign player_active = active;5�_�   L   N           M   <       ����                                                                                                                                                                                                                                                                                                                                                             d
MI     �   ;   =   ?      ) assign player_column = sprite_column_ff;5�_�   M   O           N   ;       ����                                                                                                                                                                                                                                                                                                                                                             d
MJ     �   :   <   ?      # assign player_row = sprite_row_ff;5�_�   N   P           O   :       ����                                                                                                                                                                                                                                                                                                                                                             d
MK     �   9   ;   ?      ' assign player_output = player_pix_reg;5�_�   O   Q           P   9       ����                                                                                                                                                                                                                                                                                                                                                             d
ML     �   8   :   ?       end  5�_�   P   R           Q   8       ����                                                                                                                                                                                                                                                                                                                                                             d
MO     �   7   9   ?           end5�_�   Q   S           R   7       ����                                                                                                                                                                                                                                                                                                                                                             d
MQ     �   6   8   ?      &         player_pix_reg <= player_pix;5�_�   R   T           S   6       ����                                                                                                                                                                                                                                                                                                                                                             d
MR     �   5   7   ?      +         sprite_column_ff <= btn_column_ff;5�_�   S   U           T   5       ����                                                                                                                                                                                                                                                                                                                                                             d
MR     �   4   6   ?      %         sprite_row_ff <= btn_row_ff;5�_�   T   V           U   4       ����                                                                                                                                                                                                                                                                                                                                                             d
MS     �   3   5   ?      %         btn_column_ff <= btn_column;5�_�   U   W           V   3       ����                                                                                                                                                                                                                                                                                                                                                             d
MT     �   2   4   ?              btn_row_ff <= btn_row;5�_�   V   X           W   +       ����                                                                                                                                                                                                                                                                                                                                                             d
Md     �   *   +                  btn_row_ff <= 0;5�_�   W   Y           X   +       ����                                                                                                                                                                                                                                                                                                                                                             d
Me     �   *   +                  btn_column_ff <= 0;5�_�   X   Z           Y   1       ����                                                                                                                                                                                                                                                                                                                                                             d
Mg     �   0   1                  btn_row_ff <= btn_row;5�_�   Y   [           Z   1       ����                                                                                                                                                                                                                                                                                                                                                             d
Mh    �   0   1          $        btn_column_ff <= btn_column;5�_�   Z   \           [   6        ����                                                                                                                                                                                                                                                                                                                                                             d
OS     �   5   9   ;      &assign player_output = player_pix_reg;5�_�   [   ]           \   7        ����                                                                                                                                                                                                                                                                                                                                                             d
OV     �   6   :   =       5�_�   \   ^           ]   8       ����                                                                                                                                                                                                                                                                                                                                                             d
OY     �   6   9   ?      & 83 assign sprite_row = sprite_row_ff;   (assign sprite_column = sprite_column_ff;�   7   9   ?      , 84 assign sprite_column = sprite_column_ff;5�_�   ]   _           ^   7       ����                                                                                                                                                                                                                                                                                                                                                             d
O\     �   6   8   ?      & 83 assign sprite_row = sprite_row_ff;5�_�   ^   `           _   8       ����                                                                                                                                                                                                                                                                                                                                                             d
O^     �   7   9   ?      ) assign sprite_column = sprite_column_ff;5�_�   _   a           `   ?        ����                                                                                                                                                                                                                                                                                                                                                             d
Ob     �   >               5�_�   `   b           a   9        ����                                                                                                                                                                                                                                                                                                                                                             d
Og     �   7   9   ?      (assign sprite_column = sprite_column_ff;    �   8   :   ?       5�_�   a   c           b   9       ����                                                                                                                                                                                                                                                                                                                                                             d
O�     �   8   :   >      &assign player_output = player_pix_reg;5�_�   b   d           c   9       ����                                                                                                                                                                                                                                                                                                                                                             d
O�     �   8   :   >      &assign player_output = alien2_pix_reg;5�_�   c   e           d   :       ����                                                                                                                                                                                                                                                                                                                                                             d
O�     �   9   ;   >      "assign player_row = sprite_row_ff;5�_�   d   f           e   :       ����                                                                                                                                                                                                                                                                                                                                                             d
O�     �   9   ;   >      !assign alien_row = sprite_row_ff;5�_�   e   g           f   ;       ����                                                                                                                                                                                                                                                                                                                                                             d
O�     �   :   <   >      (assign player_column = sprite_column_ff;5�_�   f   h           g   <       ����                                                                                                                                                                                                                                                                                                                                                             d
O�     �   ;   =   >      assign player_active = active;5�_�   g   i           h          ����                                                                                                                                                                                                                                                                                                                                                             d
O�    �   
      >      -    output logic   [11:0]      alien2_column,5�_�   h   j           i   
       ����                                                                                                                                                                                                                                                                                                                                                             d
QC     �   	      >      *    output logic   [11:0]      alien2_row,5�_�   i   k           j   
       ����                                                                                                                                                                                                                                                                                                                                                             d
QF     �   	      ?          5�_�   j   l           k      )    ����                                                                                                                                                                                                                                                                                                                                                             d
Qe     �   
      ?      *    output logic   [11:0]      alien2_row,�         ?    5�_�   k   m           l          ����                                                                                                                                                                                                                                                                                                                                                             d
Qk     �   
      ?      +    output logic   [11:0]      alien2_row,a   alien2_column,�         ?      -    output logic   [11:0]      alien2_column,5�_�   l   n           m   
       ����                                                                                                                                                                                                                                                                                                                                                             d
Qz     �   	      >      (    input  logic               pix_row, 5�_�   m   o           n   
   %    ����                                                                                                                                                                                                                                                                                                                                                             d
Q    �   	      >      .    input  logic   [11:0]            pix_row, 5�_�   n   p           o           ����                                                                                                                                                                                                                                                                                                                                                             d
U�    �                logic   [5:0]       counter;5�_�   o   q           p           ����                                                                                                                                                                                                                                                                                                                                                             d
V\     �      =   =       �          =    5�_�   p   r           q           ����                                                                                                                                                                                                                                                                                                                                                             d
V^     �                always_comb begin5�_�   q   s           r   
   "    ����                                                                                                                                                                                                                                                                                                                                                             d
Vo     �   	      Y      (    input  logic   [11:0]      pix_row, 5�_�   r   t           s   
   )    ����                                                                                                                                                                                                                                                                                                                                                             d
Vr     �   	      Y      *    input  logic   [11:0]      pixel_row, 5�_�   s   u           t           ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �                :// Counter for pixel number: 8x8 Grid for Alien_2 = 64 pix5�_�   t   w           u          ����                                                                                                                                                                                                                                                                                                                                                             d
V�    �         X      #logic   [11:0]      alien2_row_reg;5�_�   u   x   v       w           ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �      (   X      logic   [11:0]      _row_reg;�         X    5�_�   w   y           x           ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         n      ,l    logic   [11:0]              sprite_row;5�_�   x   |           y          ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �                +    logic   [11:0]              btn_row_ff;5�_�   y   ~   z       |          ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �                .    logic   [11:0]              btn_column_ff;5�_�   |      }       ~           ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         l      /    logic   [3:0]               player_pix_reg;5�_�   ~   �                      ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         l      .    logic   [3:0]               layer_pix_reg;5�_�      �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         l      -    logic   [3:0]               ayer_pix_reg;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         l      ,    logic   [3:0]               yer_pix_reg;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         l      +    logic   [3:0]               er_pix_reg;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         l      *    logic   [3:0]               r_pix_reg;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         l      )    logic   [3:0]               _pix_reg;5�_�   �   �           �      &    ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         l      +    logic   [3:0]               player_pix;5�_�   �   �           �      &    ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         l      1    logic                       player_active_ff;5�_�   �   �           �      
    ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         l          player_active_ff = 1'b0;5�_�   �   �           �      
    ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         l          player_pix = 4'b0000;5�_�   �   �           �      
    ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         l          player_pix_reg = 4'b0000;5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                                                             d
W     �       !              btn_column_ff = 0;5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                                                             d
W     �       !              btn_row_ff = 0;5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                                                             d
W
     �   "   #          ogic   [11:0]      _row_reg;5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                                                             d
W     �   "   #          &logic   [11:0]      alien2_column_reg;5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                                                             d
W     �   "   #          logic               active;5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                                                             d
W     �   "   #           5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                                                             d
W     �   "   #           5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                                                             d
W     �   "   #           5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                                                             d
W     �   "   #           5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                                                             d
W     �   "   #          initial begin5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                                                             d
W     �   "   #          active = 1'b0;5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                                                             d
W     �   "   #          end5�_�   �   �           �   #        ����                                                                                                                                                                                                                                                                                                                                                             d
W     �   "   #               5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      +    logic   [11:0]              sprite_row;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      *   logic   [11:0]              sprite_row;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      )  logic   [11:0]              sprite_row;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      ( logic   [11:0]              sprite_row;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      .    logic   [11:0]              sprite_column;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      -   logic   [11:0]              sprite_column;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      ,  logic   [11:0]              sprite_column;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      + logic   [11:0]              sprite_column;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      .    logic   [11:0]              sprite_row_ff;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      -   logic   [11:0]              sprite_row_ff;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      ,  logic   [11:0]              sprite_row_ff;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      + logic   [11:0]              sprite_row_ff;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      1    logic   [11:0]              sprite_column_ff;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      0   logic   [11:0]              sprite_column_ff;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      /  logic   [11:0]              sprite_column_ff;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      . logic   [11:0]              sprite_column_ff;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      /    logic   [3:0]               alien2_pix_reg;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      .   logic   [3:0]               alien2_pix_reg;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      -  logic   [3:0]               alien2_pix_reg;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      , logic   [3:0]               alien2_pix_reg;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      +    logic   [3:0]               alien2_pix;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      *   logic   [3:0]               alien2_pix;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      )  logic   [3:0]               alien2_pix;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      ( logic   [3:0]               alien2_pix;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      1    logic                       alien2_active_ff;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      0   logic                       alien2_active_ff;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      /  logic                       alien2_active_ff;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      . logic                       alien2_active_ff;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      '    logic                       active;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      &   logic                       active;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      %  logic                       active;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W     �         ^      $ logic                       active;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W      �         ^          initial begin5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W      �         ^         initial begin5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W!     �         ^        initial begin5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
W!     �         ^       initial begin5�_�   �   �           �   !        ����                                                                                                                                                                                                                                                                                                                                                             d
W$     �       "   ^          end5�_�   �   �           �   !        ����                                                                                                                                                                                                                                                                                                                                                             d
W$     �       "   ^         end5�_�   �   �           �   !        ����                                                                                                                                                                                                                                                                                                                                                             d
W$     �       "   ^        end5�_�   �   �           �   !        ����                                                                                                                                                                                                                                                                                                                                                             d
W$     �       "   ^       end5�_�   �   �           �   '        ����                                                                                                                                                                                                                                                                                                                                                             d
WM     �   R   T          %        player_pix_reg <= player_pix;�   L   N                  player_pix_reg <= 0;�   =   ?          !            player_pix = 4'b0000;�   8   :          !            player_pix = 4'b1111;�   2   4          !            player_pix = 4'b1111;�   ,   .          !            player_pix = 4'b1111;�   &   (          !            player_pix = 4'b1111;5�_�   �   �           �   S   $    ����                                                                                                                                                                                                                                                                                                                                                             d
Wn     �   R   T   ^      %        alien2_pix_reg <= player_pix;5�_�   �   �           �   R   *    ����                                                                                                                                                                                                                                                                                                                                                             d
W�     �   O   Q   ]      	    begin    �   P   R   ^      $        sprite_row_ff <= btn_row_ff;    �   Q   S   ^      *        sprite_column_ff <= btn_column_ff;5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                                                             d
W�     �   J   K                  sprite_row_ff <= 0;5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                                                             d
W�     �   J   K                  sprite_column_ff <= 0;5�_�   �   �           �   O       ����                                                                                                                                                                                                                                                                                                                                                             d
W�     �   O   Q   Z    �   O   P   Z    5�_�   �   �           �   P        ����                                                                                                                                                                                                                                                                                                                                                             d
W�     �   O   Q   [      assign alien2_active = active;5�_�   �   �           �   P        ����                                                                                                                                                                                                                                                                                                                                                             d
W�     �   O   Q   [      alien2_active = active;5�_�   �   �           �   P       ����                                                                                                                                                                                                                                                                                                                                                             d
W�     �   O   Q   [              alien2_active = active;5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                                                             d
W�     �   K   M   [    �   K   L   [    5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                                                             d
W�    �   K   M   \               alien2_active <= active;5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
Y�     �   
             9    output logic   [11:0]      alien2_row, alien2_column,5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                             d
Y�     �         [      +logic   [3:0]               alien2_pix_reg;5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                             d
Y�     �         [      *logic   [3:0]               alien2_pix_eg;5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                             d
Y�     �         [      )logic   [3:0]               alien2_pix_g;5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                             d
Y�     �         [      (logic   [3:0]               alien2_pix_;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             d
Y�     �         [          alien2_pix_reg = 4'b0000;5�_�   �   �           �   J        ����                                                                                                                                                                                                                                                                                                                                                             d
Y�     �   U   W          &assign alien2_output = alien2_pix_reg;�   N   P          %        alien2_pix_reg <= alien2_pix;�   I   K                  alien2_pix_reg <= 0;5�_�   �   �           �   W        ����                                                                                                                                                                                                                                                                                                                                                             d
Z     �   V   W          "assign alien2_row = sprite_row_ff;5�_�   �   �           �   W        ����                                                                                                                                                                                                                                                                                                                                                             d
Z     �   V   W          (assign alien2_column = sprite_column_ff;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             d
Z3     �         Y          sprite_column_ff = 0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             d
[�     �         Y          sprite_column_ff = ;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             d
[�     �          Y          sprite_row_ff = 0;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             d
[�     �      !   Y          sprite_column_ff = 316;5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             d
[�     �      !   [          5�_�   �   �           �       5    ����                                                                                                                                                                                                                                                                                                                                                             d
[�     �      !   \      7    // and as close to center as possible Cols: 317 ,->5�_�   �   �           �       7    ����                                                                                                                                                                                                                                                                                                                                                             d
[�     �      !   \      7    // and as close to center as possible Cols: 317 <->5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
\     �      !   \      ;    // and as close to center as possible Cols: 317 <-> 3245�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             d
\
     �      !   \      8    // and close to center as possible Cols: 317 <-> 3245�_�   �   �           �       (    ����                                                                                                                                                                                                                                                                                                                                                             d
\     �      !   \      :    // and close to centered as possible Cols: 317 <-> 3245�_�   �   �           �       -    ����                                                                                                                                                                                                                                                                                                                                                             d
\     �      !   \      ;    // and close to centered as possible. Cols: 317 <-> 3245�_�   �   �           �      =    ����                                                                                                                                                                                                                                                                                                                                                             d
\     �          \      =    // Initializing Alien2 20 rows from the top of the screen5�_�   �   �           �   C        ����                                                                                                                                                                                                                                                                                                                                                             d
\I     �   @   B   [              end    �   A   C   \      e    �   B   D   \       5�_�   �   �           �   C        ����                                                                                                                                                                                                                                                                                                                                                             d
\K     �   @   B   Y              end    �   A   C   Z           �   B   D   Z       5�_�   �   �           �   &   @    ����                                                                                                                                                                                                                                                                                                                                                             d
\m     �   %   '   X      �    if (((sprite_row < pixel_row) && (pixel_row < sprite_row  + 3)) && ((sprite_column < (pixel_column + 6)) && (pixel_column < sprite_column + 8)))5�_�   �   �           �   &   @    ����                                                                                                                                                                                                                                                                                                                                                             d
\q     �   %   '   X      �    if (((sprite_row < pixel_row) && (pixel_row < sprite_row  + r23)) && ((sprite_column < (pixel_column + 6)) && (pixel_column < sprite_column + 8)))5�_�   �   �           �   &   @    ����                                                                                                                                                                                                                                                                                                                                                             d
\q     �   %   '   X      �    if (((sprite_row < pixel_row) && (pixel_row < sprite_row  + 23)) && ((sprite_column < (pixel_column + 6)) && (pixel_column < sprite_column + 8)))5�_�   �   �           �   &   @    ����                                                                                                                                                                                                                                                                                                                                                             d
\s   	 �   %   '   X      �    if (((sprite_row < pixel_row) && (pixel_row < sprite_row  + 3)) && ((sprite_column < (pixel_column + 6)) && (pixel_column < sprite_column + 8)))5�_�   �   �   �       �   &        ����                                                                                                                                                                                                                                                                                                                                                             d
_�     �   %   +   X      �    if (((sprite_row < pixel_row) && (pixel_row < sprite_row  + 2)) && ((sprite_column < (pixel_column + 6)) && (pixel_column < sprite_column + 8)))5�_�   �   �           �   &        ����                                                                                                                                                                                                                                                                                                                                                             d
_�     �   %   '   \       5�_�   �   �           �   &        ����                                                                                                                                                                                                                                                                                                                                                             d
_�     �   %   8   \       �   &   '   \    5�_�   �   �   �       �   '        ����                                                                                                                                                                                                                                                                                                                                                             d
`   
 �   &   (          9    // Player's Sprite is 10 rows by 15 columns of pixels5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                                                             d
c�     �   &   (   m      9    // Alien2's Sprite is 10 rows by 15 columns of pixels5�_�   �   �           �   '       ����                                                                                                                                                                                                                                                                                                                                                             d
c�     �   &   (   m      8    // Alien2's Sprite is 0 rows by 15 columns of pixels5�_�   �   �           �   '   $    ����                                                                                                                                                                                                                                                                                                                                                             d
c�     �   &   (   m      8    // Alien2's Sprite is 8 rows by 15 columns of pixels5�_�   �   �           �   '   $    ����                                                                                                                                                                                                                                                                                                                                                             d
c�     �   &   (   m      7    // Alien2's Sprite is 8 rows by 5 columns of pixels5�_�   �   �           �   .   >    ����                                                                                                                                                                                                                                                                                                                                                             d
d     �   -   /   m      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 15))5�_�   �   �           �   .   >    ����                                                                                                                                                                                                                                                                                                                                                             d
d     �   -   /   m      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 0) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 15))5�_�   �   �           �   .   �    ����                                                                                                                                                                                                                                                                                                                                                             d
d     �   -   /   m      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 9) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 15))5�_�   �   �           �   .   �    ����                                                                                                                                                                                                                                                                                                                                                             d
d    �   -   /   m      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 9) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 95))5�_�   �   �           �   6        ����                                                                                                                                                                                                                                                                                                                                                             d
dT     �   5   6           5�_�   �   �           �   6        ����                                                                                                                                                                                                                                                                                                                                                             d
dU     �   5   6           5�_�   �   �           �   6        ����                                                                                                                                                                                                                                                                                                                                                             d
dU     �   5   6           5�_�   �   �           �   6        ����                                                                                                                                                                                                                                                                                                                                                             d
dV     �   5   6           5�_�   �   �   �       �   7   $    ����                                                                                                                                                                                                                                                                                                                                                             d
du     �   6   8   i      �    if (((sprite_row < pixel_row) && (pixel_row < sprite_row  + 2)) && ((sprite_column < (pixel_column + 6)) && (pixel_column < sprite_column + 8)))5�_�   �   �           �   7   '    ����                                                                                                                                                                                                                                                                                                                                                             d
d}     �   6   8   i      x    if ( (pixel_row < sprite_row  + 2)) && ((sprite_column < (pixel_column + 6)) && (pixel_column < sprite_column + 8)))5�_�   �   �           �   7       ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   6   8   i      w    if ( (pixel_row < sprite_row  + 2) && ((sprite_column < (pixel_column + 6)) && (pixel_column < sprite_column + 8)))5�_�   �   �           �   7   &    ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   6   8   i      x    if ( (pixel_row == sprite_row  + 2) && ((sprite_column < (pixel_column + 6)) && (pixel_column < sprite_column + 8)))5�_�   �   �           �   6        ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   5   8   i       5�_�   �   �           �   7       ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   6   8   j              5�_�   �   �           �   8   	    ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   7   9   j      x    if ( (pixel_row == sprite_row  + 1) && ((sprite_column < (pixel_column + 6)) && (pixel_column < sprite_column + 8)))5�_�   �              �   8   +    ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   7   9   j      w    if ((pixel_row == sprite_row  + 1) && ((sprite_column < (pixel_column + 6)) && (pixel_column < sprite_column + 8)))5�_�   �                8   N    ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   7   9   j      v    if ((pixel_row == sprite_row  + 1) && (sprite_column < (pixel_column + 6)) && (pixel_column < sprite_column + 8)))5�_�                  8   L    ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   7   9   j      u    if ((pixel_row == sprite_row  + 1) && (sprite_column < (pixel_column + 3) && (pixel_column < sprite_column + 8)))5�_�                 8   8    ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   7   9   j      q    if ((pixel_row == sprite_row  + 1) && (sprite_column < (pixel_column) && (pixel_column < sprite_column + 8)))5�_�                 8   r    ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   7   9   j      u    if ((pixel_row == sprite_row  + 1) && (sprite_column + 3 < (pixel_column) && (pixel_column < sprite_column + 8)))5�_�                 8   t    ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   7   9   j      u    if ((pixel_row == sprite_row  + 1) && (sprite_column + 3 < (pixel_column) && (pixel_column < sprite_column + 6)))5�_�                 :       ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   8   :   j              begin    �   9   ;   j                  active = 1'b1;5�_�                 <       ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   ;   =   i      '    // Row three of the player's sprite5�_�                 ;       ����                                                                                                                                                                                                                                                                                                                                                             d
d�     �   :   >   i              end    5�_�    	             ?       ����                                                                                                                                                                                                                                                                                                                                                             d
e     �   >   B   k      x    else if ((sprite_row + 3 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 14))5�_�    
          	   ?       ����                                                                                                                                                                                                                                                                                                                                                             d
e	     �   >   @   m          5�_�  	            
   ?       ����                                                                                                                                                                                                                                                                                                                                                             d
e     �   ?   D   m    �   ?   @   m    5�_�  
               ?       ����                                                                                                                                                                                                                                                                                                                                                             d
e     �   >   @   q          5�_�                 ?       ����                                                                                                                                                                                                                                                                                                                                                             d
e     �   >   @   q         5�_�                 ?       ����                                                                                                                                                                                                                                                                                                                                                             d
e     �   >   @   q        5�_�                 ?        ����                                                                                                                                                                                                                                                                                                                                                             d
e     �   >   @   q       5�_�                 ?        ����                                                                                                                                                                                                                                                                                                                                                             d
e     �   >   ?           5�_�                 ?       ����                                                                                                                                                                                                                                                                                                                                                             d
e     �   >   @   p      t    if ((pixel_row == sprite_row  + 1) && (sprite_column + 3 < (pixel_column) && (pixel_column < sprite_column + 6))5�_�                 =        ����                                                                                                                                                                                                                                                                                                                                                             d
e     �   ;   =   p           �   <   >   p       5�_�                 =       ����                                                                                                                                                                                                                                                                                                                                                             d
e!     �   <   >   o      %    // Row two of the player's sprite5�_�                 =       ����                                                                                                                                                                                                                                                                                                                                                             d
e(     �   <   >   o      !    // Row two of Alien2's sprite5�_�                 >   +    ����                                                                                                                                                                                                                                                                                                                                                             d
e-     �   =   ?   o      y    else if ((pixel_row == sprite_row  + 1) && (sprite_column + 3 < (pixel_column) && (pixel_column < sprite_column + 6))5�_�                 >   A    ����                                                                                                                                                                                                                                                                                                                                                             d
eB     �   =   ?   o      y    else if ((pixel_row == sprite_row  + 2) && (sprite_column + 3 < (pixel_column) && (pixel_column < sprite_column + 6))5�_�                 >   E    ����                                                                                                                                                                                                                                                                                                                                                             d
eE     �   =   ?   o      y    else if ((pixel_row == sprite_row  + 2) && (sprite_column + 2 < (pixel_column) && (pixel_column < sprite_column + 6))5�_�                 8   @    ����                                                                                                                                                                                                                                                                                                                                                             d
eI     �   7   9   o      t    if ((pixel_row == sprite_row  + 1) && (sprite_column + 3 < (pixel_column) && (pixel_column < sprite_column + 6))5�_�                 >   v    ����                                                                                                                                                                                                                                                                                                                                                             d
eX     �   =   ?   o      x    else if ((pixel_row == sprite_row  + 2) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 6))5�_�                 <        ����                                                                                                                                                                                                                                                                                                                                                             d
eb     �   :   <   o              end       �   ;   =   o       5�_�                 @       ����                                                                                                                                                                                                                                                                                                                                                             d
ej     �   @   B   n    �   @   A   n    5�_�                 B       ����                                                                                                                                                                                                                                                                                                                                                             d
ek     �   A   B              5�_�                 A       ����                                                                                                                                                                                                                                                                                                                                                             d
en     �   @   B   n      !    // Row two of Alien2's Sprite5�_�                 B       ����                                                                                                                                                                                                                                                                                                                                                             d
e�     �   A   B          x    else if ((sprite_row + 3 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 14))5�_�                 C       ����                                                                                                                                                                                                                                                                                                                                                             d
e�     �   B   C                      active = 1'b1;5�_�    !             A       ����                                                                                                                                                                                                                                                                                                                                                             d
e�     �   A   C   l    �   A   B   l    5�_�    "         !   B   )    ����                                                                                                                                                                                                                                                                                                                                                             d
e�     �   A   C   m      x    else if ((pixel_row == sprite_row  + 2) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 7))5�_�  !  #          "   B   @    ����                                                                                                                                                                                                                                                                                                                                                             d
e�     �   A   C   m      x    else if ((pixel_row == sprite_row  + 3) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 7))5�_�  "  $          #   B   u    ����                                                                                                                                                                                                                                                                                                                                                             d
e�     �   A   C   m      x    else if ((pixel_row == sprite_row  + 3) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 7))5�_�  #  %          $   F   &    ����                                                                                                                                                                                                                                                                                                                                                             d
e�     �   E   G   m      &    // Row four of the player's sprite5�_�  $  &          %   G       ����                                                                                                                                                                                                                                                                                                                                                             d
e�     �   F   G          x    else if ((sprite_row + 4 == pixel_row) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 15))5�_�  %  '          &   F       ����                                                                                                                                                                                                                                                                                                                                                             d
e�     �   F   H   l    �   F   G   l    5�_�  &  (          '   G   )    ����                                                                                                                                                                                                                                                                                                                                                             d
e�     �   F   H   m      x    else if ((pixel_row == sprite_row  + 3) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  '  )          (   G   @    ����                                                                                                                                                                                                                                                                                                                                                             d
e�     �   F   H   m      x    else if ((pixel_row == sprite_row  + 4) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  (  *          )   G   C    ����                                                                                                                                                                                                                                                                                                                                                             d
e�     �   F   H   m      x    else if ((pixel_row == sprite_row  + 4) && (sprite_column + 333 pixel_column) && (pixel_column < sprite_column + 8))5�_�  )  +          *   G   w    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   F   H   m      y    else if ((pixel_row == sprite_row  + 4) && (sprite_column + 3 != pixel_column) && (pixel_column < sprite_column + 8))5�_�  *  ,          +   G   e    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   F   H   m      y    else if ((pixel_row == sprite_row  + 4) && (sprite_column + 3 != pixel_column) && (pixel_column < sprite_column = 6))5�_�  +  -          ,   G   v    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   F   H   m      z    else if ((pixel_row == sprite_row  + 4) && (sprite_column + 3 != pixel_column) && (pixel_column != sprite_column = 6))5�_�  ,  .          -   G   J    ����                                                                                                                                                                                                                                                                                                                                                             d
f!     �   F   H   m      z    else if ((pixel_row == sprite_row  + 4) && (sprite_column + 3 != pixel_column) && (pixel_column != sprite_column + 6))5�_�  -  /          .   G   R    ����                                                                                                                                                                                                                                                                                                                                                             d
f%     �   F   H   m      {    else if ((pixel_row == sprite_row  + 4) && (sprite_column + 3 != sprite_column) && (pixel_column != sprite_column + 6))5�_�  .  0          /   G   B    ����                                                                                                                                                                                                                                                                                                                                                             d
f)     �   F   H   m          else if ((pixel_row == sprite_row  + 4) && (sprite_column + 3 != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  /  1          0   G   6    ����                                                                                                                                                                                                                                                                                                                                                             d
f-     �   F   H   m      y    else if ((pixel_row == sprite_row  + 4) && (sprite_colum!= sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  0  2          1   G   ;    ����                                                                                                                                                                                                                                                                                                                                                             d
f3     �   F   H   m      x    else if ((pixel_row == sprite_row  + 4) && (pixel_colum!= sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  1  3          2   J       ����                                                                                                                                                                                                                                                                                                                                                             d
fB     �   I   J          !            alien2_pix = 4'b1111;5�_�  2  5          3   L       ����                                                                                                                                                                                                                                                                                                                                                             d
fL     �   K   O   l      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 11)) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 16))5�_�  3  8  4      5   K       ����                                                                                                                                                                                                                                                                                                                                                             d
fS     �   J   K          1    // Row five through 10 of the player's sprite5�_�  5  9  7      8   K       ����                                                                                                                                                                                                                                                                                                                                                             d
ff     �   K   P   m    �   K   L   m    5�_�  8  :          9   K       ����                                                                                                                                                                                                                                                                                                                                                             d
fi     �   J   K             5�_�  9  ;          :   K       ����                                                                                                                                                                                                                                                                                                                                                             d
fl     �   J   L   p      "    // Row four of Alien2's Sprite5�_�  :  t          ;   L   )    ����                                                                                                                                                                                                                                                                                                                                                             d
fr     �   K   M   p      z    else if ((pixel_row == sprite_row  + 4) && (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  ;  u  <      t   L   @    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      z    else if ((pixel_row == sprite_row  + 5) && (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  t  v          u   L   A    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      j    else if ((pixel_row == sprite_row  + 5) && (sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  u  w          v   L   a    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      u    else if ((pixel_row == sprite_row  + 5) && (sprite_column < pixel_column) && (pixel_column != sprite_column + 6))5�_�  v  x          w   L   r    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      t    else if ((pixel_row == sprite_row  + 5) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 6))5�_�  w  y          x   L   &    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      t    else if ((pixel_row == sprite_row  + 5) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 9))5�_�  x  z          y   O       ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   N   P   p         5�_�  y  {          z   P       ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   O   P          �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 11)) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 16))5�_�  z  |          {   P       ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   O   P                  begin5�_�  {  }          |   P       ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   O   P                      active = 1'b1;5�_�  |  ~          }   P       ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   O   P          !            alien2_pix = 4'b1111;5�_�  }            ~   P       ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   O   P                  end5�_�  ~  �             P       ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   O   T   k          else5�_�    �          �   P       ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   P   V   n    �   P   Q   n    5�_�  �  �          �   P       ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   O   P              5�_�  �  �  �      �   U       ����                                                                                                                                                                                                                                                                                                                                                             d
g     �   U   [   r    �   U   V   r    5�_�  �  �          �   U       ����                                                                                                                                                                                                                                                                                                                                                             d
g     �   U   [   w    �   U   V   w    5�_�  �  �          �   P       ����                                                                                                                                                                                                                                                                                                                                                             d
g     �   O   Q   |      #    // Row three of Alien2's Sprite5�_�  �  �          �   P       ����                                                                                                                                                                                                                                                                                                                                                             d
g     �   O   Q   |      "    // Row hree of Alien2's Sprite5�_�  �  �          �   P       ����                                                                                                                                                                                                                                                                                                                                                             d
g     �   O   Q   |      !    // Row ree of Alien2's Sprite5�_�  �  �          �   P       ����                                                                                                                                                                                                                                                                                                                                                             d
g     �   O   Q   |           // Row ee of Alien2's Sprite5�_�  �  �          �   P       ����                                                                                                                                                                                                                                                                                                                                                             d
g     �   O   Q   |          // Row e of Alien2's Sprite5�_�  �  �          �   P       ����                                                                                                                                                                                                                                                                                                                                                             d
g     �   O   Q   |          // Row  of Alien2's Sprite5�_�  �  �          �   Q   *    ����                                                                                                                                                                                                                                                                                                                                                             d
g!     �   P   R   |      x    else if ((pixel_row == sprite_row  + 3) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   Q   A    ����                                                                                                                                                                                                                                                                                                                                                             d
g/     �   P   R   |      x    else if ((pixel_row == sprite_row  + 6) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   Q   C    ����                                                                                                                                                                                                                                                                                                                                                             d
g3     �   P   R   |      x    else if ((pixel_row == sprite_row  + 6) && (sprite_column + 3 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   Q   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g8     �   P   R   |      y    else if ((pixel_row == sprite_row  + 6) && (sprite_column + 3 == pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   Q   V    ����                                                                                                                                                                                                                                                                                                                                                             d
g;     �   P   R   |      z    else if ((pixel_row == sprite_row  + 6) && ((sprite_column + 3 == pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   Q   g    ����                                                                                                                                                                                                                                                                                                                                                             d
gE     �   P   R   |      z    else if ((pixel_row == sprite_row  + 6) && ((sprite_column + 3 == pixel_column) || (pixel_column < sprite_column + 8))5�_�  �  �          �   Q   y    ����                                                                                                                                                                                                                                                                                                                                                             d
gS     �   P   R   |      {    else if ((pixel_row == sprite_row  + 6) && ((sprite_column + 3 == pixel_column) || (pixel_column == sprite_column + 8))5�_�  �  �          �   Q   {    ����                                                                                                                                                                                                                                                                                                                                                             d
gh     �   P   R   |      {    else if ((pixel_row == sprite_row  + 6) && ((sprite_column + 3 == pixel_column) || (pixel_column == sprite_column + 6))5�_�  �  �          �   V       ����                                                                                                                                                                                                                                                                                                                                                             d
g~     �   U   W   |      #    // Row three of Alien2's Sprite5�_�  �  �          �   W   +    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      x    else if ((pixel_row == sprite_row  + 3) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      x    else if ((pixel_row == sprite_row  + 7) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      z    else if ((pixel_row == sprite_row  + 7) && xx(sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      y    else if ((pixel_row == sprite_row  + 7) && x(sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      x    else if ((pixel_row == sprite_row  + 7) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      w    else if ((pixel_row == sprite_row  + 7) && sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      v    else if ((pixel_row == sprite_row  + 7) && prite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      u    else if ((pixel_row == sprite_row  + 7) && rite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      t    else if ((pixel_row == sprite_row  + 7) && ite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      s    else if ((pixel_row == sprite_row  + 7) && te_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      r    else if ((pixel_row == sprite_row  + 7) && e_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      q    else if ((pixel_row == sprite_row  + 7) && _column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      p    else if ((pixel_row == sprite_row  + 7) && column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      o    else if ((pixel_row == sprite_row  + 7) && olumn + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      n    else if ((pixel_row == sprite_row  + 7) && lumn + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      m    else if ((pixel_row == sprite_row  + 7) && umn + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      l    else if ((pixel_row == sprite_row  + 7) && mn + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      k    else if ((pixel_row == sprite_row  + 7) && n + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      j    else if ((pixel_row == sprite_row  + 7) &&  + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      i    else if ((pixel_row == sprite_row  + 7) && + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      h    else if ((pixel_row == sprite_row  + 7) &&  1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      g    else if ((pixel_row == sprite_row  + 7) && 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      f    else if ((pixel_row == sprite_row  + 7) &&  < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      e    else if ((pixel_row == sprite_row  + 7) && < pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      d    else if ((pixel_row == sprite_row  + 7) &&  pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      c    else if ((pixel_row == sprite_row  + 7) && pixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      b    else if ((pixel_row == sprite_row  + 7) && ixel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      a    else if ((pixel_row == sprite_row  + 7) && xel_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      `    else if ((pixel_row == sprite_row  + 7) && el_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      _    else if ((pixel_row == sprite_row  + 7) && l_column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      ^    else if ((pixel_row == sprite_row  + 7) && _column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      ]    else if ((pixel_row == sprite_row  + 7) && column) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      \    else if ((pixel_row == sprite_row  + 7) && olumn) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      [    else if ((pixel_row == sprite_row  + 7) && lumn) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      Z    else if ((pixel_row == sprite_row  + 7) && umn) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      Y    else if ((pixel_row == sprite_row  + 7) && mn) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      X    else if ((pixel_row == sprite_row  + 7) && n) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      W    else if ((pixel_row == sprite_row  + 7) && ) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      V    else if ((pixel_row == sprite_row  + 7) &&  && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      U    else if ((pixel_row == sprite_row  + 7) && && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      T    else if ((pixel_row == sprite_row  + 7) && & (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      S    else if ((pixel_row == sprite_row  + 7) &&  (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      R    else if ((pixel_row == sprite_row  + 7) && (pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      Q    else if ((pixel_row == sprite_row  + 7) && pixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      P    else if ((pixel_row == sprite_row  + 7) && ixel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      O    else if ((pixel_row == sprite_row  + 7) && xel_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      N    else if ((pixel_row == sprite_row  + 7) && el_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      M    else if ((pixel_row == sprite_row  + 7) && l_column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      L    else if ((pixel_row == sprite_row  + 7) && _column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      K    else if ((pixel_row == sprite_row  + 7) && column < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      J    else if ((pixel_row == sprite_row  + 7) && olumn < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      I    else if ((pixel_row == sprite_row  + 7) && lumn < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      H    else if ((pixel_row == sprite_row  + 7) && umn < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      G    else if ((pixel_row == sprite_row  + 7) && mn < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      F    else if ((pixel_row == sprite_row  + 7) && n < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      E    else if ((pixel_row == sprite_row  + 7) &&  < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      D    else if ((pixel_row == sprite_row  + 7) && < sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      C    else if ((pixel_row == sprite_row  + 7) &&  sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      B    else if ((pixel_row == sprite_row  + 7) && sprite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      A    else if ((pixel_row == sprite_row  + 7) && prite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      @    else if ((pixel_row == sprite_row  + 7) && rite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      ?    else if ((pixel_row == sprite_row  + 7) && ite_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      >    else if ((pixel_row == sprite_row  + 7) && te_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      =    else if ((pixel_row == sprite_row  + 7) && e_column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      <    else if ((pixel_row == sprite_row  + 7) && _column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      ;    else if ((pixel_row == sprite_row  + 7) && column + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      :    else if ((pixel_row == sprite_row  + 7) && olumn + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      9    else if ((pixel_row == sprite_row  + 7) && lumn + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      8    else if ((pixel_row == sprite_row  + 7) && umn + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      7    else if ((pixel_row == sprite_row  + 7) && mn + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      6    else if ((pixel_row == sprite_row  + 7) && n + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      5    else if ((pixel_row == sprite_row  + 7) &&  + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      4    else if ((pixel_row == sprite_row  + 7) && + 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      3    else if ((pixel_row == sprite_row  + 7) &&  8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      2    else if ((pixel_row == sprite_row  + 7) && 8))5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      1    else if ((pixel_row == sprite_row  + 7) && ))5�_�  �  �          �   W   .    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      0    else if ((pixel_row == sprite_row  + 7) && )5�_�  �  �          �   W   /    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      3    else if ((pixel_row == sprite_row  + 7) &&    )�   W   X   |    5�_�  �  �          �   W   W    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      Y    else if ((pixel_row == sprite_row  + 7) &&  (pixel_row == sprite_row  + 7) &&    )  )5�_�  �  �          �   W   R    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      T    else if ((pixel_row == sprite_row  + 7) &&  (pixel_row == sprite_row  + 7) &&  )5�_�  �  �          �   W   Q    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      T    else if ((pixel_row == sprite_row  + 7) &&  (pixel_row == sprite_row  + 7) &&  )�   W   X   |    5�_�  �  �          �   W   <    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      z    else if ((pixel_row == sprite_row  + 7) &&  (pixel_row == sprite_row  + 7) && (pixel_row == sprite_row  + 7) &&    ) )5�_�  �  �          �   W   :    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      z    else if ((pixel_row == sprite_row  + 7) &&  (pixel_row != sprite_row  + 7) && (pixel_row == sprite_row  + 7) &&    ) )5�_�  �  �          �   W   0    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      }    else if ((pixel_row == sprite_row  + 7) &&  (pixel_column != sprite_row  + 7) && (pixel_row == sprite_row  + 7) &&    ) )5�_�  �  �          �   W   ?    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      |    else if ((pixel_row == sprite_row  + 7) && (pixel_column != sprite_row  + 7) && (pixel_row == sprite_row  + 7) &&    ) )5�_�  �  �          �   W   1    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      m    else if ((pixel_row == sprite_row  + 7) && ( sprite_row  + 7) && (pixel_row == sprite_row  + 7) &&    ) )5�_�  �  �          �   W   <    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      l    else if ((pixel_row == sprite_row  + 7) && (sprite_row  + 7) && (pixel_row == sprite_row  + 7) &&    ) )5�_�  �  �          �   W   >    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      k    else if ((pixel_row == sprite_row  + 7) && (sprite_row + 7) && (pixel_row == sprite_row  + 7) &&    ) )5�_�  �  �          �   W   \    ����                                                                                                                                                                                                                                                                                                                                                             d
g�     �   V   X   |      w    else if ((pixel_row == sprite_row  + 7) && (sprite_row + 2 < pixel_row) && (pixel_row == sprite_row  + 7) &&    ) )5�_�  �  �          �   W   k    ����                                                                                                                                                                                                                                                                                                                                                             d
h      �   V   X   |      v    else if ((pixel_row == sprite_row  + 7) && (sprite_row + 2 < pixel_row) && (pixel_row < sprite_row  + 7) &&    ) )5�_�  �  �          �   W   t    ����                                                                                                                                                                                                                                                                                                                                                             d
h     �   V   X   |      u    else if ((pixel_row == sprite_row  + 7) && (sprite_row + 2 < pixel_row) && (pixel_row < sprite_row + 7) &&    ) )5�_�  �  �          �   W   t    ����                                                                                                                                                                                                                                                                                                                                                             d
h     �   V   X   |      t    else if ((pixel_row == sprite_row  + 7) && (sprite_row + 2 < pixel_row) && (pixel_row < sprite_row + 7) &&    ))5�_�  �  �          �   W   o    ����                                                                                                                                                                                                                                                                                                                                                             d
h     �   V   X   |      s    else if ((pixel_row == sprite_row  + 7) && (sprite_row + 2 < pixel_row) && (pixel_row < sprite_row + 7) &&    )5�_�  �  �          �   W   f    ����                                                                                                                                                                                                                                                                                                                                                             d
h#     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_row + 2 < pixel_row) && (pixel_row < sprite_row + 7) && (pixel_column   )5�_�  �  �          �   W   Y    ����                                                                                                                                                                                                                                                                                                                                                             d
h'     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_row + 2 < pixel_row) && (pixel_row < sprite_column + 7) && (pixel_column   )5�_�  �  �          �   W   J    ����                                                                                                                                                                                                                                                                                                                                                             d
h-     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_row + 2 < pixel_row) && (pixel_column < sprite_column + 7) && (pixel_column   )5�_�  �  �          �   W   :    ����                                                                                                                                                                                                                                                                                                                                                             d
h3     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_row + 2 < pixel_column) && (pixel_column < sprite_column + 7) && (pixel_column   )5�_�  �  �          �   W   A    ����                                                                                                                                                                                                                                                                                                                                                             d
hF     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 7) && (pixel_column   )5�_�  �  �          �   W   D    ����                                                                                                                                                                                                                                                                                                                                                             d
hX     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 7) && (pixel_column   )5�_�  �  �          �   W   B    ����                                                                                                                                                                                                                                                                                                                                                             d
h_     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_column + 1 pixel_column) && (pixel_column < sprite_column + 7) && (pixel_column   )5�_�  �  �          �   W   e    ����                                                                                                                                                                                                                                                                                                                                                             d
hk     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_column + 1 != pixel_column) && (pixel_column < sprite_column + 7) && (pixel_column   )5�_�  �  �          �   W   w    ����                                                                                                                                                                                                                                                                                                                                                             d
hr     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_column + 1 != pixel_column) && (pixel_colum != sprite_column + 7) && (pixel_column   )5�_�  �  �          �   W   b    ����                                                                                                                                                                                                                                                                                                                                                             d
hx     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_column + 1 != pixel_column) && (pixel_colum != sprite_column + 3) && (pixel_column   )5�_�  �  �          �   W   �    ����                                                                                                                                                                                                                                                                                                                                                             d
h{     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_column + 1 != pixel_column) && (pixel_column != sprite_column + 3) && (pixel_column   )5�_�  �  �          �   W   �    ����                                                                                                                                                                                                                                                                                                                                                             d
h�     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_column + 1 != pixel_column) && (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 8)   )5�_�  �  �          �   W   E    ����                                                                                                                                                                                                                                                                                                                                                             d
h�     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_column + 1 != pixel_column) && (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 8))5�_�  �  �          �   W   A    ����                                                                                                                                                                                                                                                                                                                                                             d
h�     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (sprite_column + 1pixel_column) && (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 8))5�_�  �            �   W   <    ����                                                                                                                                                                W   <                                                                                                                                                                                        d
h�     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (pixel_column) && (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 8))5�_�  �              W   J    ����                                                                                                                                                                W   <                                                                                                                                                                                        d
h�     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (pixel_column != sprite_col + 1) && (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 8))5�_�                 U       ����                                                                                                                                                                W   <                                                                                                                                                                                        d
i     �   T   U                  5�_�                 [       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i&     �   Z   [          x    else if ((pixel_row == sprite_row  + 3) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�                 Z       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i*     �   Y   \   z      #    // Row three of Alien2's Sprite5�_�                 \       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i-     �   [   ^   {              begin5�_�                 ]        ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i.     �   \   ^   |      begin5�_�    	             \       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i1     �   \   ^   |    �   \   ]   |    5�_�    
          	   \       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i4     �   [   \              5�_�  	            
   Z       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i5     �   Y   Z              5�_�  
               Z       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i<     �   Y   [   {      #    // Row three of Alien2's Sprite5�_�                 Z       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i<     �   Y   [   {      "    // Row hree of Alien2's Sprite5�_�                 Z       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i<     �   Y   [   {      !    // Row ree of Alien2's Sprite5�_�                 Z       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i<     �   Y   [   {           // Row ee of Alien2's Sprite5�_�                 Z       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i<     �   Y   [   {          // Row e of Alien2's Sprite5�_�                 Z       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i>     �   Y   [   {          // Row  of Alien2's Sprite5�_�                 [       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
iN     �   Z   [          x    else if ((pixel_row == sprite_row  + 3) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 8))5�_�                 Z       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
iS     �   Z   \   z    �   Z   [   z    5�_�                 [   )    ����                                                                                                                                                                V   <                                                                                                                                                                                        d
iW     �   Z   \   {      �    else if ((pixel_row == sprite_row  + 7) && (pixel_column != sprite_column + 1) && (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 8))5�_�                 [   P    ����                                                                                                                                                                V   <                                                                                                                                                                                        d
ij     �   Z   \   {      �    else if ((pixel_row == sprite_row  + 8) && (pixel_column != sprite_column + 1) && (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 8))5�_�                 [   w    ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i�     �   Z   \   {      �    else if ((pixel_row == sprite_row  + 8) && (pixel_column != sprite_column + 2) && (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 8))5�_�                 [   w    ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i�     �   Z   \   {      �    else if ((pixel_row == sprite_row  + 8) && (pixel_column != sprite_column + 2) && (pixel_column != sprite_column + 2) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 8))5�_�                 [   �    ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i�     �   Z   \   {      �    else if ((pixel_row == sprite_row  + 8) && (pixel_column != sprite_column + 2) && (pixel_column != sprite_column + 4) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 8))5�_�                 [   �    ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i�     �   Z   \   {      �    else if ((pixel_row == sprite_row  + 8) && (pixel_column != sprite_column + 2) && (pixel_column != sprite_column + 4) && (pixel_column != sprite_column + 5) && (pixel_column != sprite_column + 8))5�_�                 b       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i�     �   a   b                      active = 1'b0;5�_�                 _       ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i�     �   ]   _   z              end    �   ^   `   z              5�_�                 6        ����                                                                                                                                                                V   <                                                                                                                                                                                        d
i�     �   5   9   y       5�_�                 7        ����                                                                                                                                                                X   <                                                                                                                                                                                        d
i�     �   6   8   {       5�_�                 8        ����                                                                                                                                                                X   <                                                                                                                                                                                        d
i�     �   6   8   {              �   7   9   {       5�_�                        ����                                                                                                                                                                W   <                                                                                                                                                                                        d
i�     �      	   z      //5�_�                         ����                                                                                                                                                                Z   <                                                                                                                                                                                        d
i�     �         {      //    �         |      //    �         }      //    �      	   }      //5�_�    !                 0    ����                                                                                                                                                                W   <                                                                                                                                                                                        d
i�     �         z      0// Created by Alexander Maso PSU ECE-Winter 20235�_�     "          !          ����                                                                                                                                                                [   <                                                                                                                                                                                        d
i�     �      
   ~      //5�_�  !  #          "          ����                                                                                                                                                                \   <                                                                                                                                                                                        d
j     �   
            //5�_�  "              #   	       ����                                                                                                                                                                \   <                                                                                                                                                                                        d
j    �      
         // implementatio5�_�  �              W   d    ����                                                                                                                                                                                                                                                                                                                                                             d
h�     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (pixel_column != sprite_col + 1 || sprite_column + 3) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 8))5�_�                    W   D    ����                                                                                                                                                                                                                                                                                                                                                             d
h�     �   V   X   |      �    else if ((pixel_row == sprite_row  + 7) && (pixel_column != sprite_col + 1 || sprite_column + 3) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 8))5�_�  �          �  �   U       ����                                                                                                                                                                                                                                                                                                                                                             d
g     �   U   V   r    �   U   V   r          5�_�  ;  =      t  <   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f|     �   K   M   p      y    else if ((pixel_row == sprite_row  + 5) & (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  <  >          =   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      x    else if ((pixel_row == sprite_row  + 5)  (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  =  ?          >   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      w    else if ((pixel_row == sprite_row  + 5) (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  >  @          ?   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      v    else if ((pixel_row == sprite_row  + 5) pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  ?  A          @   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      u    else if ((pixel_row == sprite_row  + 5) ixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  @  B          A   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      t    else if ((pixel_row == sprite_row  + 5) xel_column != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  A  C          B   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      s    else if ((pixel_row == sprite_row  + 5) el_column != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  B  D          C   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      r    else if ((pixel_row == sprite_row  + 5) l_column != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  C  E          D   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      q    else if ((pixel_row == sprite_row  + 5) _column != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  D  F          E   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      p    else if ((pixel_row == sprite_row  + 5) column != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  E  G          F   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      o    else if ((pixel_row == sprite_row  + 5) olumn != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  F  H          G   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      n    else if ((pixel_row == sprite_row  + 5) lumn != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  G  I          H   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      m    else if ((pixel_row == sprite_row  + 5) umn != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  H  J          I   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      l    else if ((pixel_row == sprite_row  + 5) mn != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  I  K          J   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      k    else if ((pixel_row == sprite_row  + 5) n != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  J  L          K   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      j    else if ((pixel_row == sprite_row  + 5)  != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  K  M          L   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      i    else if ((pixel_row == sprite_row  + 5) != sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  L  N          M   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      h    else if ((pixel_row == sprite_row  + 5) = sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  M  O          N   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      g    else if ((pixel_row == sprite_row  + 5)  sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  N  P          O   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      f    else if ((pixel_row == sprite_row  + 5) sprite_column + 3) && (pixel_column != sprite_column + 6))5�_�  O  Q          P   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      e    else if ((pixel_row == sprite_row  + 5) prite_column + 3) && (pixel_column != sprite_column + 6))5�_�  P  R          Q   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      d    else if ((pixel_row == sprite_row  + 5) rite_column + 3) && (pixel_column != sprite_column + 6))5�_�  Q  S          R   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      c    else if ((pixel_row == sprite_row  + 5) ite_column + 3) && (pixel_column != sprite_column + 6))5�_�  R  T          S   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      b    else if ((pixel_row == sprite_row  + 5) te_column + 3) && (pixel_column != sprite_column + 6))5�_�  S  U          T   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      a    else if ((pixel_row == sprite_row  + 5) e_column + 3) && (pixel_column != sprite_column + 6))5�_�  T  V          U   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f}     �   K   M   p      `    else if ((pixel_row == sprite_row  + 5) _column + 3) && (pixel_column != sprite_column + 6))5�_�  U  W          V   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      _    else if ((pixel_row == sprite_row  + 5) column + 3) && (pixel_column != sprite_column + 6))5�_�  V  X          W   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      ^    else if ((pixel_row == sprite_row  + 5) olumn + 3) && (pixel_column != sprite_column + 6))5�_�  W  Y          X   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      ]    else if ((pixel_row == sprite_row  + 5) lumn + 3) && (pixel_column != sprite_column + 6))5�_�  X  Z          Y   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      \    else if ((pixel_row == sprite_row  + 5) umn + 3) && (pixel_column != sprite_column + 6))5�_�  Y  [          Z   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      [    else if ((pixel_row == sprite_row  + 5) mn + 3) && (pixel_column != sprite_column + 6))5�_�  Z  \          [   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      Z    else if ((pixel_row == sprite_row  + 5) n + 3) && (pixel_column != sprite_column + 6))5�_�  [  ]          \   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      Y    else if ((pixel_row == sprite_row  + 5)  + 3) && (pixel_column != sprite_column + 6))5�_�  \  ^          ]   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      X    else if ((pixel_row == sprite_row  + 5) + 3) && (pixel_column != sprite_column + 6))5�_�  ]  _          ^   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      W    else if ((pixel_row == sprite_row  + 5)  3) && (pixel_column != sprite_column + 6))5�_�  ^  `          _   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      V    else if ((pixel_row == sprite_row  + 5) 3) && (pixel_column != sprite_column + 6))5�_�  _  a          `   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      U    else if ((pixel_row == sprite_row  + 5) ) && (pixel_column != sprite_column + 6))5�_�  `  b          a   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      T    else if ((pixel_row == sprite_row  + 5)  && (pixel_column != sprite_column + 6))5�_�  a  c          b   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      S    else if ((pixel_row == sprite_row  + 5) && (pixel_column != sprite_column + 6))5�_�  b  d          c   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      R    else if ((pixel_row == sprite_row  + 5) & (pixel_column != sprite_column + 6))5�_�  c  e          d   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f     �   K   M   p      Q    else if ((pixel_row == sprite_row  + 5)  (pixel_column != sprite_column + 6))5�_�  d  f          e   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      P    else if ((pixel_row == sprite_row  + 5) (pixel_column != sprite_column + 6))5�_�  e  g          f   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      O    else if ((pixel_row == sprite_row  + 5) pixel_column != sprite_column + 6))5�_�  f  h          g   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      N    else if ((pixel_row == sprite_row  + 5) ixel_column != sprite_column + 6))5�_�  g  i          h   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      M    else if ((pixel_row == sprite_row  + 5) xel_column != sprite_column + 6))5�_�  h  j          i   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      L    else if ((pixel_row == sprite_row  + 5) el_column != sprite_column + 6))5�_�  i  k          j   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      K    else if ((pixel_row == sprite_row  + 5) l_column != sprite_column + 6))5�_�  j  l          k   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      J    else if ((pixel_row == sprite_row  + 5) _column != sprite_column + 6))5�_�  k  m          l   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      I    else if ((pixel_row == sprite_row  + 5) column != sprite_column + 6))5�_�  l  n          m   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      H    else if ((pixel_row == sprite_row  + 5) olumn != sprite_column + 6))5�_�  m  o          n   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      G    else if ((pixel_row == sprite_row  + 5) lumn != sprite_column + 6))5�_�  n  p          o   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      F    else if ((pixel_row == sprite_row  + 5) umn != sprite_column + 6))5�_�  o  q          p   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      E    else if ((pixel_row == sprite_row  + 5) mn != sprite_column + 6))5�_�  p  r          q   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      D    else if ((pixel_row == sprite_row  + 5) n != sprite_column + 6))5�_�  q  s          r   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      C    else if ((pixel_row == sprite_row  + 5)  != sprite_column + 6))5�_�  r              s   L   ,    ����                                                                                                                                                                                                                                                                                                                                                             d
f�     �   K   M   p      B    else if ((pixel_row == sprite_row  + 5) != sprite_column + 6))5�_�  5      6  8  7   K       ����                                                                                                                                                                                                                                                                                                                                                             d
fX     �   K   L   m    �   K   L   m      1    // Row five through 10 of the player's sprite5�_�  5          7  6   J       ����                                                                                                                                                                                                                                                                                                                                                             d
fT     �   J   K   m    �   J   K   m      1    // Row five through 10 of the player's sprite5�_�  3          5  4   K       ����                                                                                                                                                                                                                                                                                                                                                             d
fO     �   K   L   n    �   K   L   n      "    // Row four of Alien2's Sprite   z    else if ((pixel_row == sprite_row  + 4) && (pixel_column != sprite_column + 3) && (pixel_column != sprite_column + 6))           begin               active = 1'b1;5�_�            !      B   )    ����                                                                                                                                                                                                                                                                                                                                                             d
e�     �   A   C   m      x    else if ((pixel_row == sprite_row  + 3) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 7))5�_�   �           �   �   6        ����                                                                                                                                                                                                                                                                                                                                                             d
dY     �   5   8        5�_�   �           �   �   '        ����                                                                                                                                                                                                                                                                                                                                                             d
`
     �   &   (          9    // Alien2's Sprite is 10 rows by 15 columns of pixels5�_�   �           �   �   %        ����                                                                                                                                                                                                                                                                                                                                                             d
_�     �   %   &   X    �   $   &   X      Fa    // Enable output of the player's sprite when in the proper region   9    // Player's Sprite is 10 rows by 15 columns of pixels   G    // *** Still unsure on the implementation of this active signal....   P    // ...Do I want to just use two assignments with a ternary operator instead?       //    :    // assign active = (sprite_row < pixel row) && .......   4    // assign player_active = active ? 1'b1 : 1'b0;        //   �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 15))           begin               active = 1'b1;           end       else           begin               active = 1'b0;           end       lways_comb begin5�_�   |           ~   }           ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         l      !    logic   [3:0]               ;5�_�   y   {       |   z          ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �              5�_�   z               {          ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �              5�_�   u           w   v           ����                                                                                                                                                                                                                                                                                                                                                             d
V�     �         X    �         X      ,/    logic   [11:0]              sprite_row;   .    logic   [11:0]              sprite_column;   .    logic   [11:0]              sprite_row_ff;   1    logic   [11:0]              sprite_column_ff;   +    logic   [11:0]              btn_row_ff;   .    logic   [11:0]              btn_column_ff;   /    logic   [3:0]               player_pix_reg;   +    logic   [3:0]               player_pix;   1    logic                       player_active_ff;   '    logic                       active;              initial begin       active = 1'b0;       player_active_ff = 1'b0;       player_pix = 4'b0000;       player_pix_reg = 4'b0000;       sprite_column_ff = 0;       sprite_row_ff = 0;       btn_column_ff = 0;       btn_row_ff = 0;       end       / Internals5��