Vim�UnDo� �	����VfcW�E�]��N�C]�^΄d��89   �       player_row = 431;   !         v       v   v   v    d�`    _�                     '       ����                                                                                                                                                                                                                                                                                                                                                             d��     �   &   '          <    // Alien2's Sprite is 16 rows by 16 columns of pixels   5�_�                       H    ����                                                                                                                                                                                                                                                                                                                                                             d�     �          �      R    // Initializing Player 20 rows from the bottom of the screen. Rows 451 <-> 4605�_�                       H    ����                                                                                                                                                                                                                                                                                                                                                             d�
     �          �      N    // Initializing Player 20 rows from the bottom of the screen. Rows 4-> 4605�_�                       K    ����                                                                                                                                                                                                                                                                                                                                                             d�     �          �      R    // Initializing Player 20 rows from the bottom of the screen. Rows 441 --> 4605�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d�     �          �      S    // Initializing Player 20 rows from the bottom of the screen. Rows 441 <--> 4605�_�                       I    ����                                                                                                                                                                                                                                                                                                                                                             d�      �          �      S    // Initializing Player 30 rows from the bottom of the screen. Rows 441 <--> 4605�_�                       R    ����                                                                                                                                                                                                                                                                                                                                                             d�"     �          �      S    // Initializing Player 30 rows from the bottom of the screen. Rows 431 <--> 4605�_�      	              '       ����                                                                                                                                                                                                                                                                                                                                                             d�5     �   &   (   �         5�_�      
           	   '   /    ����                                                                                                                                                                                                                                                                                                                                                             d�V     �   &   (   �      6    // Player sprite is 20 rows by 30 columns (pixels)5�_�   	              
   )       ����                                                                                                                                                                                                                                                                                                                                                             d�`     �   (   )          J    // ***** TURN THIS INTO AN ASSIGN STATEMEN WITH TERNARY OPERATOR *****5�_�   
                 )   O    ����                                                                                                                                                                                                                                                                                                                                                             d�g     �   (   *   �      �    player_active_reg = ((player_row < pixel_row) && (pixel_row < player_row + 11) && (player_column < pixel_column) && (pixel_column < player_column + 16));5�_�                    )   �    ����                                                                                                                                                                                                                                                                                                                                                             d�q     �   (   *   �      �    player_active_reg = ((player_row < pixel_row) && (pixel_row < player_row + 21) && (player_column < pixel_column) && (pixel_column < player_column + 16));5�_�                    )   �    ����                                                                                                                                                                                                                                                                                                                                                             d�r     �   (   *   �      �    player_active_reg = ((player_row < pixel_row) && (pixel_row < player_row + 21) && (player_column < pixel_column) && (pixel_column < player_column + 6));5�_�                    )   �    ����                                                                                                                                                                                                                                                                                                                                                             d�s     �   (   *   �      �    player_active_reg = ((player_row < pixel_row) && (pixel_row < player_row + 21) && (player_column < pixel_column) && (pixel_column < player_column + ));5�_�                    -       ����                                                                                                                                                                                                                                                                                                                                                             d�	     �   ,   .   �      9    // Row one and two of the player's sprite            5�_�                   .   ?    ����                                                                                                                                                                                                                                                                                                                                                             d�.     �   -   /   �      i    if ((player_row < pixel_row) && (pixel_row < player_row  + 3) && (pixel_column == player_column + 8))5�_�                    .   h    ����                                                                                                                                                                                                                                                                                                                            .   E       .   g       v   g    d�8     �   -   /   �      i    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column == player_column + 8))�   .   /   �    5�_�                    .   h    ����                                                                                                                                                                                                                                                                                                                            .   E       .   g       v   g    d�=     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column == player_column + 8))(pixel_column == player_column + 8)5�_�                    .   h    ����                                                                                                                                                                                                                                                                                                                            .   E       .   g       v   g    d�>     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column == player_column + 8)(pixel_column == player_column + 8)5�_�                    .   |    ����                                                                                                                                                                                                                                                                                                                            .   E       .   g       v   g    d�A     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column == player_column + 8) && (pixel_column == player_column + 8)5�_�                    .   �    ����                                                                                                                                                                                                                                                                                                                            .   E       .   g       v   g    d�I     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column == player_column + 8) && (pixel_column < player_column + 8)5�_�                    .   �    ����                                                                                                                                                                                                                                                                                                                            .   E       .   g       v   g    d�X     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column == player_column + 8) && (pixel_column < player_column + 17)5�_�                    .   U    ����                                                                                                                                                                                                                                                                                                                            .   E       .   g       v   g    d�^     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column == player_column + 8) && (pixel_column < player_column + 17))5�_�                    .   f    ����                                                                                                                                                                                                                                                                                                                            .   E       .   g       v   g    d�c     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < player_column + 8) && (pixel_column < player_column + 17))5�_�                    .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�u     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < player_column + 14) && (pixel_column < player_column + 17))5�_�                    .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < layer_column + 14) && (pixel_column < player_column + 17))5�_�                    .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < ayer_column + 14) && (pixel_column < player_column + 17))5�_�                    .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < yer_column + 14) && (pixel_column < player_column + 17))5�_�                     .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < er_column + 14) && (pixel_column < player_column + 17))5�_�      !               .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < r_column + 14) && (pixel_column < player_column + 17))5�_�       "           !   .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < _column + 14) && (pixel_column < player_column + 17))5�_�   !   #           "   .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < column + 14) && (pixel_column < player_column + 17))5�_�   "   $           #   .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < olumn + 14) && (pixel_column < player_column + 17))5�_�   #   %           $   .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < lumn + 14) && (pixel_column < player_column + 17))5�_�   $   &           %   .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < umn + 14) && (pixel_column < player_column + 17))5�_�   %   '           &   .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < mn + 14) && (pixel_column < player_column + 17))5�_�   &   (           '   .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < n + 14) && (pixel_column < player_column + 17))5�_�   '   )           (   .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column <  + 14) && (pixel_column < player_column + 17))5�_�   (   *           )   .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < + 14) && (pixel_column < player_column + 17))5�_�   )   +           *   .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column <  14) && (pixel_column < player_column + 17))5�_�   *   2           +   .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < 14) && (pixel_column < player_column + 17))5�_�   +   3   1       2   .   V    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dǊ     �   -   /   �          if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < 4) && (pixel_column < player_column + 17))5�_�   2   4           3   .   F    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dǎ     �   -   /   �      {    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column) && (pixel_column < player_column + 17))5�_�   3   5           4   2       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dǱ     �   1   3   �      '    // Row three of the player's sprite5�_�   4   6           5   2       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d��     �   2   4   �    �   2   3   �    5�_�   5   7           6   3       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d��     �   2   4   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (player_column + 14 < pixel_column) && (pixel_column < player_column + 17))5�_�   6   8           7   3       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d��     �   2   4   �      �    else if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (player_column + 14 < pixel_column) && (pixel_column < player_column + 17))5�_�   7   9           8   2       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�     �   1   3   �      (    // Rows 3 & 4 of the player's sprite5�_�   8   :           9   2       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�     �   1   3   �      (    // Rows 3 & 6 of the player's sprite5�_�   9   ;           :   3       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�     �   2   4   �      �    else if ((player_row + 2 < pixel_row) && (pixel_row < player_row  + 5) && (player_column + 14 < pixel_column) && (pixel_column < player_column + 17))5�_�   :   <           ;   3   J    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�     �   2   4   �      �    else if ((player_row + 4 < pixel_row) && (pixel_row < player_row  + 5) && (player_column + 14 < pixel_column) && (pixel_column < player_column + 17))5�_�   ;   =           <   3   `    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�     �   2   4   �      �    else if ((player_row + 4 < pixel_row) && (pixel_row < player_row  + 7) && (player_column + 14 < pixel_column) && (pixel_column < player_column + 17))5�_�   <   >           =   3   �    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�M     �   2   4   �      �    else if ((player_row + 4 < pixel_row) && (pixel_row < player_row  + 7) && (player_column + 4 < pixel_column) && (pixel_column < player_column + 17))5�_�   =   ?           >   4       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�Q     �   3   4          x    else if ((player_row + 3 == pixel_row) && (player_column + 2 < pixel_column) && (pixel_column < player_column + 14))5�_�   >   @           ?   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �      &    // Row four of the player's sprite5�_�   ?   A           @   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �      %    // Row our of the player's sprite5�_�   @   B           A   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �      $    // Row ur of the player's sprite5�_�   A   C           B   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �      #    // Row r of the player's sprite5�_�   B   D           C   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �      "    // Row  of the player's sprite5�_�   C   E           D   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �      !    // Row of the player's sprite5�_�   D   F           E   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �           // Row f the player's sprite5�_�   E   G           F   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �          // Row  the player's sprite5�_�   F   H           G   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �          // Row the player's sprite5�_�   G   I           H   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �          // Row he player's sprite5�_�   H   J           I   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �          // Row e player's sprite5�_�   I   K           J   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �          // Row  player's sprite5�_�   J   L           K   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �          // Row player's sprite5�_�   K   M           L   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�`     �   6   8   �          // Row layer's sprite5�_�   L   N           M   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�a     �   6   8   �          // Row ayer's sprite5�_�   M   O           N   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�a     �   6   8   �          // Row yer's sprite5�_�   N   P           O   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�a     �   6   8   �          // Row er's sprite5�_�   O   Q           P   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�a     �   6   8   �          // Row r's sprite5�_�   P   R           Q   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�a     �   6   8   �          // Row 's sprite5�_�   Q   S           R   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�b     �   6   8   �          // Row s sprite5�_�   R   T           S   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�b     �   6   8   �          // Row  sprite5�_�   S   U           T   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�b     �   6   8   �          // Row sprite5�_�   T   V           U   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�b     �   6   8   �          // Row prite5�_�   U   W           V   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�b     �   6   8   �          // Row rite5�_�   V   X           W   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�b     �   6   8   �          // Row ite5�_�   W   Y           X   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�b     �   6   8   �          // Row te5�_�   X   Z           Y   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�b     �   6   8   �          // Row e5�_�   Y   [           Z   7   
    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�c     �   6   8   �          // Row �   7   8   �    5�_�   Z   \           [   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�e     �   6   8   �          // Row e5�_�   [   ]           \   7   
    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�i     �   7   9   �    �   7   8   �    5�_�   \   ^           ]   7   
    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�m     �   6   8   �          // Row 5�_�   ]   _           ^   7       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�q     �   6   8   �          // Rows 5�_�   ^   `           _   9       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�}     �   8   9          x    else if ((player_row + 4 == pixel_row) && (player_column + 1 < pixel_column) && (pixel_column < player_column + 15))5�_�   _   a           `   8       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dȃ     �   7   9   �      �    else if ((player_row + 4 < pixel_row) && (pixel_row < player_row  + 7) && (player_column + 4 < pixel_column) && (pixel_column < player_column + 27))5�_�   `   b           a   8   J    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dȇ     �   7   9   �      �    else if ((player_row + 6 < pixel_row) && (pixel_row < player_row  + 7) && (player_column + 4 < pixel_column) && (pixel_column < player_column + 27))5�_�   a   c           b   8   `    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dȐ     �   7   9   �      �    else if ((player_row + 6 < pixel_row) && (pixel_row < player_row  + 9) && (player_column + 4 < pixel_column) && (pixel_column < player_column + 27))5�_�   b   d           c   8   �    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dȗ     �   7   9   �      �    else if ((player_row + 6 < pixel_row) && (pixel_row < player_row  + 9) && (player_column + 2 < pixel_column) && (pixel_column < player_column + 27))5�_�   c   e           d   <        ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dȫ     �   <   ?   �    �   <   =   �    5�_�   d   f           e   <       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dȮ     �   ;   <          1    // Row five through 10 of the player's sprite5�_�   e   h           f   >       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dȱ     �   =   >          �    else if (((player_row + 4 < pixel_row) && (pixel_row < player_row  + 11)) && (player_column < pixel_column) && (pixel_column < player_column + 16))5�_�   f   i   g       h   <       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dȹ     �   ;   =   �          // Rows 7 & 85�_�   h   j           i   <       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dȼ     �   ;   =   �          // Rows 9 & 85�_�   i   k           j   <       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d��     �   ;   =   �          // Rows 9 & 15�_�   j   l           k   =       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d��     �   <   >   �      �    else if ((player_row + 6 < pixel_row) && (pixel_row < player_row  + 9) && (player_column + 2 < pixel_column) && (pixel_column < player_column + 29))5�_�   k   m           l   =   I    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d��     �   <   >   �      �    else if ((player_row + 8 < pixel_row) && (pixel_row < player_row  + 9) && (player_column + 2 < pixel_column) && (pixel_column < player_column + 29))5�_�   l   n           m   <       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d��     �   ;   =   �          // Rows 9 & 105�_�   m   o           n   <       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d��     �   ;   =   �          // Rows 9 -205�_�   n   p           o   =   I    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d��     �   <   >   �      �    else if ((player_row + 8 < pixel_row) && (pixel_row < player_row  + 11) && (player_column + 2 < pixel_column) && (pixel_column < player_column + 29))5�_�   o   q           p   =   a    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d��     �   <   >   �      �    else if ((player_row + 8 < pixel_row) && (pixel_row < player_row  + 21) && (player_column + 2 < pixel_column) && (pixel_column < player_column + 29))5�_�   p   r           q   =   �    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d��     �   <   >   �      �    else if ((player_row + 8 < pixel_row) && (pixel_row < player_row  + 21) && (player_column < pixel_column) && (pixel_column < player_column + 29))5�_�   q   s           r   !       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�      �       "   �          player_row = 460;5�_�   r   t           s       6    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�F     �      !   �      >    // and close to centered as possible. Columns: 313 <-> 3285�_�   s   u           t       >    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�K     �      !   �      >    // and close to centered as possible. Columns: 306 <-> 3285�_�   t   v           u   "       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�W     �   !   #   �          player_column = 312;5�_�   u               v   !       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�_    �       "   �          player_row = 431;5�_�   f           h   g   =       ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dȳ     �   <   ?        5�_�   +       ,   2   1   .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    dǅ     �   .   /   �    �   -   /   �      �    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < 4 ) && (pixel_column < player_column + 17))5�_�   +   -       1   ,   .   U    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�v     �   -   /   �      ~    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column < ) && (pixel_column < player_column + 17))5�_�   ,   .           -   .   S    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�w     �   -   /   �      }    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column  ) && (pixel_column < player_column + 17))5�_�   -   /           .   .   R    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�x     �   -   /   �      |    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column ) && (pixel_column < player_column + 17))5�_�   .   0           /   .   R    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�z     �   -   /   �      {    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column) && (pixel_column < player_column + 17))5�_�   /               0   .   F    ����                                                                                                                                                                                                                                                                                                                            .   U       .   f       v   f    d�|     �   .   /   �    �   -   /   �      |    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (p ixel_column) && (pixel_column < player_column + 17))5�_�                   .   @    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   -   /   �      i    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && (pixel_column == player_column + 8))5�_�                     .   U    ����                                                                                                                                                                                                                                                                                                                                                             d�%     �   -   /   �      Z    if ((player_row < pixel_row) && (pixel_row < player_row  + 5) && ( player_column + 8))5��