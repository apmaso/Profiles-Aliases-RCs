Vim�UnDo� ��&��09��#�)�����p�����>�   v   �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 15))   5   ?      �       �   �   �    d
d;    _�                             ����                                                                                                                                                                                                                                                                                                                                                             d
N     �   0   2          �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < ship_row + 11)) && (sprite_column < pixel_column) && (pixel_column < ship_column + 16))�                 �    if (((sprite_row < pixel_row) && (pixel_row < ship_row + 3)) && ((sprite_column < (pixel_column + 6)) && (pixel_column < ship_column + 8)))5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d
N8     �   0   2          �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 11)) && (sprite_column < pixel_column) && (pixel_column < ship_column + 16))�   *   ,          v    else if ((sprite_row + 4 == pixel_row) && (sprite_column + 1 < pixel_column) && (pixel_column < ship_column + 15))�   $   &          v    else if ((sprite_row + 3 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < ship_column + 14))�                 �    if (((sprite_row < pixel_row) && (pixel_row < sprite_row  + 3)) && ((sprite_column < (pixel_column + 6)) && (pixel_column < ship_column + 8)))5�_�                          ����                                                                                                                                                                                                                                                                                                                                                             d
N�     �         V    �         V    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
N�     �                1    logic   [11:0]              sprite_column_ff;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
N�     �         W    �         W    5�_�                       -    ����                                                                                                                                                                                                                                                                                                                                                             d
N�     �         X      .    logic   [11:0]              sprite_row_ff;5�_�      	                 0    ����                                                                                                                                                                                                                                                                                                                                                             d
N�     �         X      1    logic   [11:0]              sprite_column_ff;5�_�      
           	   V       ����                                                                                                                                                                                                                                                                                                                                                             d
N�     �   U   W   X      assign player_active = active;5�_�   	              
   R        ����                                                                                                                                                                                                                                                                                                                                                             d
N�     �   R   T   X    �   R   S   X    5�_�   
                 R        ����                                                                                                                                                                                                                                                                                                                                                             d
N�     �   R   T   Y    �   R   S   Y    5�_�                    S       ����                                                                                                                                                                                                                                                                                                                                                             d
N�     �   R   T   Z      "assign player_row = sprite_row_ff;5�_�                    T       ����                                                                                                                                                                                                                                                                                                                                                             d
N�    �   S   U   Z      (assign player_column = sprite_column_ff;5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             d
R�     �   	      Z      :    output logic [11:0]         player_row, player_column,5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             d
R�     �   	      Z      3    logic [11:0]         player_row, player_column,5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             d
R�     �   	      Z      9    input logic [11:0]         player_row, player_column,5�_�                    
   &    ����                                                                                                                                                                                                                                                                                                                                                             d
R�     �   	      Z      :    input logic  [11:0]         player_row, player_column,5�_�                    
   1    ����                                                                                                                                                                                                                                                                                                                                                             d
R�     �   	      Z      9    input logic  [11:0]         pixel_row, player_column,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
S+     �         Z    �         Z    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d
S7     �         [      '    logic                       active;5�_�                       -    ����                                                                                                                                                                                                                                                                                                                                                             d
S:     �         [      .    logic                       player_active;5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                             d
SB     �         [    �         [    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
SD     �                1    logic                       player_active_ff;5�_�                    Y       ����                                                                                                                                                                                                                                                                                                                                                             d
SY     �   X   Z   [      assign player_active = active;5�_�                    Y   $    ����                                                                                                                                                                                                                                                                                                                                                             d
S^     �   X   Z   [      %assign player_active = player_active;5�_�                    P   %    ����                                                                                                                                                                                                                                                                                                                                                             d
Sb     �   O   R   [      %        player_pix_reg <= player_pix;5�_�                    H       ����                                                                                                                                                                                                                                                                                                                                                             d
S�     �   H   J   \    �   H   I   \    5�_�                    I       ����                                                                                                                                                                                                                                                                                                                                                             d
S�     �   H   J   ]      #        player_active_ff <= active;5�_�                    I       ����                                                                                                                                                                                                                                                                                                                                                             d
S�    �   H   J   ]              player_active_ff <= ;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
T     �         ]          end5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d
T     �         ^          5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                             d
T*     �         ^          player_pix = 4'b0000;5�_�       "           !          ����                                                                                                                                                                                                                                                                                                                                                             d
T/     �         _    �         _    5�_�   !   #           "           ����                                                                                                                                                                                                                                                                                                                                                             d
T1     �                 5�_�   "   $           #          ����                                                                                                                                                                                                                                                                                                                                                             d
T4     �         _          player_pix = 4'b0000;5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                                             d
TF     �         _    �         _    5�_�   $   &           %          ����                                                                                                                                                                                                                                                                                                                                                             d
TJ     �         `          player_pix_reg = 4'b0000;5�_�   %   '           &          ����                                                                                                                                                                                                                                                                                                                                                             d
T\     �         `          player_active_ff = 4'b0000;5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                                             d
T_     �         `          player_active_ff = 1'b0000;5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                             d
T~     �         `      1    logic   [11:0]              sprite_column_ff;5�_�   (   *           )          ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �         `      0    logic   [11:0]             sprite_column_ff;5�_�   )   ,           *          ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �      !   `          player_pix_reg = 4'b0000;5�_�   *   -   +       ,            ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �      !   a       �       !   a    5�_�   ,   .           -            ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �      !   a      sprite_column_ff5�_�   -   /           .            ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �      !   a      sprite_column_ff5�_�   .   0           /           ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �      "   a          sprite_column_ff5�_�   /   1           0   !        ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �   !   #   b    �   !   "   b    5�_�   0   2           1   !        ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �       !           5�_�   1   3           2   !       ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �       "   b          sprite_column_ff = 0;5�_�   2   4           3   !       ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �       "   b          sprite_= 0;5�_�   3   5           4   !       ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �       "   b          sprite_row_ff= 0;5�_�   4   6           5   !       ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �   !   %   b    �   !   "   b    5�_�   5   7           6   $       ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �   #   $              end5�_�   6   8           7   "   
    ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �   !   #   d          sprite_column_ff = 0;5�_�   7   =           8   #   
    ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �   "   $   d          sprite_row_ff = 0;5�_�   8   >   ;       =          ����                                                                                                                                                                                                                                                                                                                                                             d
U?     �         d      //5�_�   =   @           >          ����                                                                                                                                                                                                                                                                                                                                                             d
U@     �         f      //5�_�   >   A   ?       @      )    ����                                                                                                                                                                                                                                                                                                                                                             d
V     �         h      *// asynchronous for the different sprites?5�_�   @   C           A      *    ����                                                                                                                                                                                                                                                                                                                                                             d
V    �         h      *// asynchronous for the different sprites?5�_�   A   D   B       C           ����                                                                                                                                                                                                                                                                                                                                                             d
YJ    �   b   d          &assign player_output = player_pix_reg;�   [   ]          %        player_pix_reg <= player_pix;�   R   T                  player_pix_reg <= 0;�   "   $              player_pix_reg = 4'b0000;�                /    logic   [3:0]               player_pix_reg;5�_�   C   E           D   -   l    ����                                                                                                                                                                                                                                                                                                                                                             d
\�     �   ,   .   h      �    if (((sprite_row < pixel_row) && (pixel_row < sprite_row  + 3)) && ((sprite_column < (pixel_column + 6)) && (pixel_column < sprite_column + 8)))5�_�   D   F           E   -   V    ����                                                                                                                                                                                                                                                                                                                                                             d
\�     �   ,   .   h      k    if (((sprite_row < pixel_row) && (pixel_row < sprite_row  + 3)) && (pixel_column < sprite_column + 8)))5�_�   E   G           F   3   .    ����                                                                                                                                                                                                                                                                                                                                                             d
\�     �   2   4   h      x    else if ((sprite_row + 3 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 14))5�_�   F   H           G   3   /    ����                                                                                                                                                                                                                                                                                                                                                             d
\�     �   2   4   h      y    else if ((sprite_row + 3 == pixel_row) && ((sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 14))5�_�   G   I           H   -   C    ����                                                                                                                                                                                                                                                                                                                                                             d
\�     �   ,   .   h      l    if (((sprite_row < pixel_row) && (pixel_row < sprite_row  + 3)) && (pixel_column == sprite_column + 8)))5�_�   H   J           I   -   
    ����                                                                                                                                                                                                                                                                                                                                                             d
\�     �   ,   .   h      k    if (((sprite_row < pixel_row) && (pixel_row < sprite_row  + 3) && (pixel_column == sprite_column + 8)))5�_�   I   K           J   /       ����                                                                                                                                                                                                                                                                                                                                                             d
]6     �   .   /                      active = 1'b1;5�_�   J   L           K   4       ����                                                                                                                                                                                                                                                                                                                                                             d
]8     �   3   4                      active = 1'b1;5�_�   K   M           L   9       ����                                                                                                                                                                                                                                                                                                                                                             d
]9     �   8   9                      active = 1'b1;5�_�   L   N           M   >       ����                                                                                                                                                                                                                                                                                                                                                             d
];     �   =   >                      active = 1'b1;5�_�   M   O           N   B       ����                                                                                                                                                                                                                                                                                                                                                             d
]<     �   A   B                      active = 1'b0;5�_�   N   P           O   ,       ����                                                                                                                                                                                                                                                                                                                                                             d
]B     �   +   /   c          always_comb begin5�_�   O   Q           P   -        ����                                                                                                                                                                                                                                                                                                                                                             d
]E     �   ,   /   e       5�_�   P   R           Q   .   #    ����                                                                                                                                                                                                                                                                                                                                                             d
]�     �   -   /   f      $    if ((sprite_row < pixel_row) && 5�_�   Q   S           R   .   F    ����                                                                                                                                                                                                                                                                                                                                                             d
]�     �   -   /   f      S    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (pixel_column 5�_�   R   T           S   .   b    ����                                                                                                                                                                                                                                                                                                                                                             d
]�     �   -   /   f      c    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (sprite_column < pixel_column 5�_�   S   U           T   .   B    ����                                                                                                                                                                                                                                                                                                                                                             d
]�     �   -   /   f      d    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (sprite_column < pixel_column) 5�_�   T   V           U   .   c    ����                                                                                                                                                                                                                                                                                                                                                             d
]�     �   -   /   f      d    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (sprite_column < pixel_column) �   .   /   f    5�_�   U   W           V   .   e    ����                                                                                                                                                                                                                                                                                                                                                             d
]�     �   -   /   f      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (sprite_column < pixel_column)  && (sprite_column < pixel_column) 5�_�   V   X           W   .   n    ����                                                                                                                                                                                                                                                                                                                                                             d
]�     �   -   /   f      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (sprite_column < pixel_column) && (sprite_column < pixel_column) 5�_�   W   Y           X   .   |    ����                                                                                                                                                                                                                                                                                                                                                             d
]�     �   -   /   f      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (sprite_column < pixel_column) && (pixel_column < pixel_column) 5�_�   X   Z           Y   .   �    ����                                                                                                                                                                                                                                                                                                                                                             d
]�     �   -   /   f      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (sprite_column < pixel_column) && (pixel_column < sprite_column) 5�_�   Y   [           Z   .   �    ����                                                                                                                                                                                                                                                                                                                                                             d
]�     �   -   0   f      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 15) 5�_�   Z   \           [   -   E    ����                                                                                                                                                                                                                                                                                                                                                             d
^     �   ,   /   g      E    // Enable output of the player's sprite when in the proper region5�_�   [   ]           \   .   9    ����                                                                                                                                                                                                                                                                                                                                                             d
^!     �   -   0   h      9    // Player's Sprite is 10 rows by 15 columns of pixels5�_�   \   ^           ]   /       ����                                                                                                                                                                                                                                                                                                                                                             d
^%     �   -   /   i      9    // Player's Sprite is 10 rows by 15 columns of pixels    �   .   0   i          //5�_�   ]   _           ^   0       ����                                                                                                                                                                                                                                                                                                                                                             d
^*     �   /   3   h             active = 0 5�_�   ^   `           _   0       ����                                                                                                                                                                                                                                                                                                                                                             d
^4     �   /   1   j             active = 0;5�_�   _   a           `   1       ����                                                                                                                                                                                                                                                                                                                                                             d
^5     �   0   2   j          else5�_�   `   b           a   0       ����                                                                                                                                                                                                                                                                                                                                                             d
^<     �   /   2   j             active = 0;5�_�   a   c           b   0       ����                                                                                                                                                                                                                                                                                                                                                             d
^?     �   /   1   k          5�_�   b   d           c   1       ����                                                                                                                                                                                                                                                                                                                                                             d
^D     �   0   2   k              active = 0;5�_�   c   e           d   1       ����                                                                                                                                                                                                                                                                                                                                                             d
^G     �   0   3   k                  active = 0;5�_�   d   f           e   3       ����                                                                                                                                                                                                                                                                                                                                                             d
^K     �   2   6   l          else5�_�   e   g           f   4       ����                                                                                                                                                                                                                                                                                                                                                             d
^R     �   3   5   n      	    begin5�_�   f   h           g   5       ����                                                                                                                                                                                                                                                                                                                                                             d
^S     �   4   6   n              5�_�   g   i           h   1       ����                                                                                                                                                                                                                                                                                                                                                             d
^]     �   0   2   n                  active = 0;5�_�   h   j           i   5       ����                                                                                                                                                                                                                                                                                                                                                             d
^d     �   4   8   n                  active = 1'b0;5�_�   i   k           j   /       ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   .   1   p      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 15))5�_�   j   l           k   /       ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   .   1   q          5�_�   k   m           l   0   !    ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   /   1   r      O    // ......Do I want to just us an assignment and a ternary operator instead?5�_�   l   n           m   0   %    ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   /   1   r      P    // ......Do I want to just use an assignment and a ternary operator instead?5�_�   m   o           n   0   1    ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   /   1   r      Q    // ......Do I want to just use two assignment and a ternary operator instead?5�_�   n   p           o   0   6    ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   /   1   r      R    // ......Do I want to just use two assignments and a ternary operator instead?5�_�   o   q           p   0   S    ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   /   4   r      S    // ......Do I want to just use two assignments with a ternary operator instead?5�_�   p   r           q   2       ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   1   3   u          //5�_�   q   s           r   1       ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   0   2   u          //5�_�   r   t           s   0   
    ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   /   1   u      S    // ......Do I want to just use two assignments with a ternary operator instead?5�_�   s   u           t   1       ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   0   3   u          //  5�_�   t   v           u   2       ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   1   3   v      !    // active_bool = (sprite_row 5�_�   u   w           v   2       ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   1   3   v          // active_bool = (�   2   3   v    5�_�   v   x           w   2        ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   1   3   v      !    // active_bool = (sprite_row �   2   3   v    5�_�   w   y           x   2   !    ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   1   3   v      ,    // active_bool = (sprite_row sprite_row 5�_�   x   z           y   2        ����                                                                                                                                                                                                                                                                                                                                                             d
^�     �   1   3   v      !    // active_bool = (sprite_row 5�_�   y   {           z   2   8    ����                                                                                                                                                                                                                                                                                                                                                             d
_
     �   1   4   v      9    // active_bool = (sprite_row < pixel row) && ....... 5�_�   z   |           {   4       ����                                                                                                                                                                                                                                                                                                                                                             d
_     �   2   4   w          //    �   3   5   w          //  5�_�   {   }           |   2       ����                                                                                                                                                                                                                                                                                                                                                             d
_     �   1   3   v      8    // active_bool = (sprite_row < pixel row) && .......5�_�   |   ~           }   2       ����                                                                                                                                                                                                                                                                                                                                                             d
_$     �   1   3   v      ?    // assign active_bool = (sprite_row < pixel row) && .......5�_�   }              ~   3       ����                                                                                                                                                                                                                                                                                                                                                             d
_(     �   2   4   v          // assign aci 5�_�   ~   �              3       ����                                                                                                                                                                                                                                                                                                                                                             d
_*     �   2   4   v          // assign player_aci 5�_�      �           �   3       ����                                                                                                                                                                                                                                                                                                                                                             d
_+    �   2   4   v          // assign player_acti 5�_�   �   �           �   5   ?    ����                                                                                                                                                                                                                                                                                                                                                             d
d"     �   4   6   v      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 10) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 15))5�_�   �               �   5   �    ����                                                                                                                                                                                                                                                                                                                                                             d
d:    �   4   6   v      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 11) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 15))5�_�   A           C   B   ,       ����                                                                                                                                                                                                                                                                                                                            ,          ,          v        d
V%     �   +   L   h      ,    always_ff @ (posedge clk or posedge rst)�   +   -   I      -    ualways_ff @ (posedge clk or posedge rst)5�_�   >           @   ?      *    ����                                                                                                                                                                                                                                                                                                                                                             d
U�    �         h      /// asynchronous for the different sprites?  ***5�_�   8   <   9   =   ;          ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �              5�_�   ;               <          ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �              5�_�   8   :       ;   9          ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �              5�_�   9               :          ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �              5�_�   *           ,   +          ����                                                                                                                                                                                                                                                                                                                                                             d
T�     �          a    �          a      -    psprite_column_fflayer_pix_reg = 4'b0000;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
N�     �         V    �         V      .    logic   [11:0]              sprite_row_ff;   1    logic   [11:0]              sprite_column_ff;5��