Vim�UnDo� Wι��}��>�B�n��=��i��M2��6�E�   V                  x       x   x   x    d
J�    _�                             ����                                                                                                                                                                                                                                                                                                                                                             d
=a     �                   5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d
=j     �       	         D    // ship is centered in the upper left corner | Row x Col / (0,0)5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d
=~    �      	   !      A:// ship is centered in the upper left corner | Row x Col / (0,0)5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d
A     �          !       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
AI     �         "      // in my SpaceInvaders5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d
AL     �         "      // in my Space Invaders5�_�                       <    ����                                                                                                                                                                                                                                                                                                                                                             d
A^     �          "      <// SystemVerilog Module for the "Earth Defender" (or Player)5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             d
Ak     �         "      // in t Space Invaders5�_�      
           	           ����                                                                                                                                                                                                                                                                                                                                                            d
A�     �      	   %       5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                            d
A�     �      
   &      module 5�_�   
                    !    ����                                                                                                                                                                                                                                                                                                                                                            d
B[     �      
   (      !    input logic         clk, rst,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            d
B     �      	   )      (    input logic         clk, rst, enable5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                            d
B�     �      
   )          output logic [11:0]5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            d
B�     �      	   )      -    input logic              clk, rst, enable5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                            d
B�     �         )          output logic [11:0]     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                            d
B�     �   
      +      )5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            d
B�     �   
      +          )5�_�                            ����                                                                                                                                                                                                                                                                                                                                                            d
C�     �   #   %          �    else if (((ship_row + 4 < pixel_row) && (pixel_row < ship_row + 11)) && (ship_column < pixel_column) && (pixel_column < ship_column + 16))�                 r    else if ((ship_row + 4 == pixel_row) && (ship_column + 1 < pixel_column) && (pixel_column < ship_column + 15))�                r    else if ((ship_row + 3 == pixel_row) && (ship_column + 2 < pixel_column) && (pixel_column < ship_column + 14))�                �    if (((ship_row < pixel_row) && (pixel_row < ship_row + 3)) && ((ship_column < (pixel_column + 6)) && (pixel_column < ship_column + 8)))5�_�                            ����                                                                                                                                                                                                                                                                                                                                                            d
D     �   #   %          �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < ship_row + 11)) && (ship_column < pixel_column) && (pixel_column < ship_column + 16))�                 t    else if ((sprite_row + 4 == pixel_row) && (ship_column + 1 < pixel_column) && (pixel_column < ship_column + 15))�                t    else if ((sprite_row + 3 == pixel_row) && (ship_column + 2 < pixel_column) && (pixel_column < ship_column + 14))�                �    if (((sprite_row < pixel_row) && (pixel_row < ship_row + 3)) && ((ship_column < (pixel_column + 6)) && (pixel_column < ship_column + 8)))5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            d
D     �                    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                            d
D     �         *      @// ship is centered in the upper left corner | Row x Col / (0,0)5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            d
D     �         *          5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                            d
D;     �         +    �         +    5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                            d
D?     �         ,      +    logic   [11:0]              sprite_row;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                            d
Ds     �   *   ,          !            vga_output = 4'b0000;�   &   (          !            vga_output = 4'b1111;�   !   #          !            vga_output = 4'b1111;�                !            vga_output = 4'b1111;�                !            vga_output = 4'b1111;5�_�                    ,       ����                                                                                                                                                                                                                                                                                                                                                            d
D�     �   +                  end5�_�                    -        ����                                                                                                                                                                                                                                                                                                                                                            d
D�     �   ,   0   /       5�_�                    /        ����                                                                                                                                                                                                                                                                                                                                                            d
D�     �   .   <   1       5�_�                            ����                                                                                                                                                                                                                                                                                                                                                            d
D�     �         =       5�_�                    /       ����                                                                                                                                                                                                                                                                                                                                                            d
D�     �   .   0   =      7always_ff @ (posedge vga_fast_clk or posedge vga_rst_i)5�_�                     =        ����                                                                                                                                                                                                                                                                                                                                                            d
D�     �   <               5�_�      !                  0    ����                                                                                                                                                                                                                                                                                                                                                            d
D�     �      
   =      0    input logic                 clk, rst, enable5�_�       "           !          ����                                                                                                                                                                                                                                                                                                                                                            d
E     �         >    �         >    5�_�   !   #           "           ����                                                                                                                                                                                                                                                                                                                                                            d
E     �         @      +    logic   [11:0]              sprite_row;5�_�   "   $           #           ����                                                                                                                                                                                                                                                                                                                                                            d
E      �         @      !    logic   [11:0]              ;5�_�   #   %           $      -    ����                                                                                                                                                                                                                                                                                                                                                            d
E.     �         @      .    logic   [11:0]              sprite_column;5�_�   $   &           %   	   0    ����                                                                                                                                                                                                                                                                                                                                                            d
E8     �      
   @      0    input logic  [11:0]         btn_row, btn_col5�_�   %   '           &   <       ����                                                                                                                                                                                                                                                                                                                                                            d
EE     �   ;   =   @              btn_col_ff <= btn_col;5�_�   &   (           '   <       ����                                                                                                                                                                                                                                                                                                                                                            d
EI     �   ;   =   @      !        btn_col_ff <= btn_column;5�_�   '   )           (   7       ����                                                                                                                                                                                                                                                                                                                                                            d
EO     �   6   8   @              btn_col_ff <= 0;5�_�   (   *           )   7       ����                                                                                                                                                                                                                                                                                                                                                            d
EP     �   6   8   @              btn_col_ff <= 0;5�_�   )   +           *   4       ����                                                                                                                                                                                                                                                                                                                                                            d
EX     �   3   5   @          if (vga_rst_i)5�_�   *   ,           +   4       ����                                                                                                                                                                                                                                                                                                                                                            d
E[     �   3   5   @          if (rst_i)5�_�   +   -           ,   2       ����                                                                                                                                                                                                                                                                                                                                                            d
E^     �   1   3   @      always_ff @ (posedge5�_�   ,   .           -   ?        ����                                                                                                                                                                                                                                                                                                                                                            d
Ej     �   >   B   @       5�_�   -   /           .   @        ����                                                                                                                                                                                                                                                                                                                                                            d
Em     �   >   @   B           �   ?   A   B       5�_�   .   0           /      *    ����                                                                                                                                                                                                                                                                                                                                                            d
E�     �         A      +    logic   [11:0]              sprite_row;5�_�   /   1           0      -    ����                                                                                                                                                                                                                                                                                                                                                            d
E�     �         A      .    logic   [11:0]              sprite_column;5�_�   0   2           1   ;       ����                                                                                                                                                                                                                                                                                                                                                            d
E�     �   ;   >   A    �   ;   <   A    5�_�   1   3           2   =       ����                                                                                                                                                                                                                                                                                                                                                            d
E�     �   <   >   C      $        btn_column_ff <= btn_column;5�_�   2   4           3   =       ����                                                                                                                                                                                                                                                                                                                                                            d
E�     �   <   >   C      #        btn_olumn_ff <= btn_column;5�_�   3   5           4   =       ����                                                                                                                                                                                                                                                                                                                                                            d
E�     �   <   >   C              btn_<= btn_column;5�_�   4   6           5   =       ����                                                                                                                                                                                                                                                                                                                                                            d
E�     �   <   >   C               btn_row_ff<= btn_column;5�_�   5   7           6   <       ����                                                                                                                                                                                                                                                                                                                                                            d
E�     �   ;   =   C              btn_row_ff <= btn_row;5�_�   6   8           7   <        ����                                                                                                                                                                                                                                                                                                                                                            d
E�     �   ;   =   C      !        btn_column_ff <= btn_row;5�_�   7   9           8   <       ����                                                                                                                                                                                                                                                                                                                                                            d
E�     �   ;   =   C      '        btn_column_ff <= btn_column_ff;5�_�   8   :           9   ;       ����                                                                                                                                                                                                                                                                                                                                                            d
E�     �   :   <   C              btn_row_ff <= btn_row;5�_�   9   ;           :   ;       ����                                                                                                                                                                                                                                                                                                                                                            d
E�     �   :   <   C      !        btn_row_ff <= btn_row_ff;5�_�   :   <           ;          ����                                                                                                                                                                                                                                                                                                                                                            d
F3     �         C    �         C    5�_�   ;   =           <          ����                                                                                                                                                                                                                                                                                                                                                            d
F5     �                    always_comb begin5�_�   <   >           =          ����                                                                                                                                                                                                                                                                                                                                                            d
F8     �         C      D    // ship is centered in the upper left corner | Row x Col / (0,0)5�_�   =   ?           >          ����                                                                                                                                                                                                                                                                                                                                                            d
F?     �         C      #    // Row three of the ship sprite5�_�   >   @           ?   "       ����                                                                                                                                                                                                                                                                                                                                                            d
FD     �   !   #   C      "    // Row four of the ship sprite5�_�   ?   A           @   '   '    ����                                                                                                                                                                                                                                                                                                                                                            d
FL     �   &   (   C      -    // Row five through 10 of the ship sprite5�_�   @   B           A      0    ����                                                                                                                                                                                                                                                                                                                                                            d
G�     �      	   C      0    input logic                 clk, rst, enable5�_�   A   C           B      *    ����                                                                                                                                                                                                                                                                                                                                                            d
G�     �   
      C      *    output logic [3:0]          player_pix5�_�   B   D           C           ����                                                                                                                                                                                                                                                                                                                                                            d
G�     �         C       5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                                                            d
G�     �         C    �         C    5�_�   D   F           E          ����                                                                                                                                                                                                                                                                                                                                                            d
G�     �         D      -    output logic [3:0]          player_output5�_�   E   G           F      	    ����                                                                                                                                                                                                                                                                                                                                                            d
G�     �         D      &    logic [3:0]          player_output5�_�   F   H           G          ����                                                                                                                                                                                                                                                                                                                                                            d
G�     �         D      )    logic    [3:0]          player_output5�_�   G   I           H          ����                                                                                                                                                                                                                                                                                                                                                            d
G�     �         D      (    logic   [3:0]          player_output5�_�   H   J           I      -    ����                                                                                                                                                                                                                                                                                                                                                            d
G�     �         D      -    logic   [3:0]               player_output5�_�   I   K           J      *    ����                                                                                                                                                                                                                                                                                                                                                            d
G�     �         D      -    logic   [3:0]               player_pixff;5�_�   J   L           K          ����                                                                                                                                                                                                                                                                                                                                                            d
H!     �         D    �         D    5�_�   K   M           L          ����                                                                                                                                                                                                                                                                                                                                                            d
H#     �                    5�_�   L   N           M      -    ����                                                                                                                                                                                                                                                                                                                                                            d
H'     �         D      .    logic   [3:0]               player_pix_ff;5�_�   M   O           N      -    ����                                                                                                                                                                                                                                                                                                                                                            d
H>     �         D      .    logic   [3:0]               player_pix_ff;5�_�   N   P           O   ?       ����                                                                                                                                                                                                                                                                                                                                                            d
HW     �   ?   B   D    �   ?   @   D    5�_�   O   Q           P   <       ����                                                                                                                                                                                                                                                                                                                                                            d
HY     �   ;   <          $        sprite_row_ff <= btn_row_ff;5�_�   P   S           Q   <       ����                                                                                                                                                                                                                                                                                                                                                            d
HZ     �   ;   <          *        sprite_column_ff <= btn_column_ff;5�_�   Q   T   R       S   <       ����                                                                                                                                                                                                                                                                                                                                                            d
Ho     �   ;   =   D              btn_row_ff<= btn_row;5�_�   S   U           T   @       ����                                                                                                                                                                                                                                                                                                                                                            d
Hw     �   ?   B   D              end5�_�   T   V           U   A       ����                                                                                                                                                                                                                                                                                                                                                            d
H{     �   @   B   E          end5�_�   U   W           V   @       ����                                                                                                                                                                                                                                                                                                                                                            d
H�     �   ?   A   E              5�_�   V   X           W   8       ����                                                                                                                                                                                                                                                                                                                                                            d
H�     �   8   <   E    �   8   9   E    5�_�   W   Y           X   9       ����                                                                                                                                                                                                                                                                                                                                                            d
H�     �   8   :   H      $        sprite_row_ff <= btn_row_ff;5�_�   X   Z           Y   :       ����                                                                                                                                                                                                                                                                                                                                                            d
H�     �   9   ;   H      *        sprite_column_ff <= btn_column_ff;5�_�   Y   [           Z   ;       ����                                                                                                                                                                                                                                                                                                                                                            d
H�     �   :   <   H      %        player_pix_reg <= player_pix;5�_�   Z   \           [   ;       ����                                                                                                                                                                                                                                                                                                                                                            d
H�     �   :   <   H              player_pix_reg <= ;5�_�   [   ]           \   :       ����                                                                                                                                                                                                                                                                                                                                                            d
H�     �   9   ;   H              sprite_column_ff <= ;5�_�   \   ^           ]   9       ����                                                                                                                                                                                                                                                                                                                                                            d
H�     �   8   :   H              sprite_row_ff <= ;5�_�   ]   _           ^   G        ����                                                                                                                                                                                                                                                                                                                                                            d
H�     �   F   I   H       5�_�   ^   `           _   G       ����                                                                                                                                                                                                                                                                                                                                                            d
H�     �   F   H   I      a5�_�   _   a           `   G       ����                                                                                                                                                                                                                                                                                                                                                            d
H�     �   F   H   I      assign 5�_�   `   b           a   G   &    ����                                                                                                                                                                                                                                                                                                                                                            d
I	     �   F   I   I      &assign player_output = player_pix_reg;5�_�   a   c           b   H   !    ����                                                                                                                                                                                                                                                                                                                                                            d
I     �   H   J   J    �   H   I   J    5�_�   b   d           c   I       ����                                                                                                                                                                                                                                                                                                                                                            d
I!     �   H   J   K      "assign player_row = sprite_row_ff;5�_�   c   e           d   I   !    ����                                                                                                                                                                                                                                                                                                                                                            d
I&     �   H   J   K      %assign player_column = sprite_row_ff;5�_�   d   f           e   
   6    ����                                                                                                                                                                                                                                                                                                                                                            d
I6     �   	      K      7    output logic [11:0]         player_row, player_col,5�_�   e   g           f      -    ����                                                                                                                                                                                                                                                                                                                                                            d
I?     �   
      K      -    output logic [3:0]          player_output5�_�   f   h           g           ����                                                                                                                                                                                                                                                                                                                                                            d
Ie     �         L       5�_�   g   i           h           ����                                                                                                                                                                                                                                                                                                                                                            d
I�     �         M      &    output logic                active5�_�   h   j           i          ����                                                                                                                                                                                                                                                                                                                                                            d
I�     �         M          5�_�   i   k           j          ����                                                                                                                                                                                                                                                                                                                                                            d
I�     �         M              begin5�_�   j   l           k           ����                                                                                                                                                                                                                                                                                                                                                            d
I�     �         N       5�_�   k   m           l           ����                                                                                                                                                                                                                                                                                                                                                            d
I�     �      !   P                  active = 1'b1;5�_�   l   n           m   %       ����                                                                                                                                                                                                                                                                                                                                                            d
I�     �   %   '   P    �   %   &   P    5�_�   m   o           n   +       ����                                                                                                                                                                                                                                                                                                                                                            d
I�     �   +   -   Q    �   +   ,   Q    5�_�   n   p           o   1       ����                                                                                                                                                                                                                                                                                                                                                            d
I�     �   1   3   R    �   1   2   R    5�_�   o   q           p   6       ����                                                                                                                                                                                                                                                                                                                                                            d
I�     �   6   8   S    �   6   7   S    5�_�   p   s           q   9       ����                                                                                                                                                                                                                                                                                                                                                            d
I�     �   8   :   T          end5�_�   q   t   r       s   7       ����                                                                                                                                                                                                                                                                                                                                                            d
I�     �   6   8   T                  active = 1'b1;5�_�   s   u           t   S        ����                                                                                                                                                                                                                                                                                                                                                            d
Jk     �   R   U   T       5�_�   t   v           u   S        ����                                                                                                                                                                                                                                                                                                                                                            d
Jl     �   R   T   U       5�_�   u   w           v          ����                                                                                                                                                                                                                                                                                                                                                            d
J�     �         U              active = 1'b0;5�_�   v   x           w          ����                                                                                                                                                                                                                                                                                                                                                            d
J�     �         U              active = 1'b0;5�_�   w               x           ����                                                                                                                                                                                                                                                                                                                                                            d
J�    �         U       5�_�   q           s   r   7       ����                                                                                                                                                                                                                                                                                                                                                            d
I�     �   6   8   T                  active = 1'01;5�_�   Q           S   R   8       ����                                                                                                                                                                                                                                                                                                                                                            d
H^     �   8   9   D    �   8   9   D      *        sprite_column_ff <= btn_column_ff;5��