Vim�UnDo� /Ψ3�{&��W
�4#�9a���c��A���    ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 42 == pixel_column) || (sprite_column + 45 == pixel_column) || (pixel_column == sprite_column + 46) || (pixel_column == sprite_column + 51) || (pixel_column == sprite_column + 52)))   �  =      N       N   N   N    d�]    _�                     T   H    ����                                                                                                                                                                                                                                                                                                                                                             d�E     �   S   U       7    else if ((sprite_row + 6 < pixel_row) && (pixel_row < sprite_row  +  9) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 5)) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 12 < pixel_column) && (pixel_column < sprite_column + 17))))5�_�                    T   D    ����                                                                                                                                                                                                                                                                                                                                                             d�G     �   S   U       6    else if ((sprite_row + 6 < pixel_row) && (pixel_row < sprite_row  + 9) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 5)) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 12 < pixel_column) && (pixel_column < sprite_column + 17))))5�_�                    c   b    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   b   d       <    else if ((sprite_row + 12 < pixel_row) && (pixel_row < sprite_row  + 15) && ((sprite_column + 2 == pixel_column) || (sprite_column + 3 == pixel_column) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    c   �    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   b   d       <    else if ((sprite_row + 12 < pixel_row) && (pixel_row < sprite_row  + 15) && ((sprite_column + 3 == pixel_column) || (sprite_column + 3 == pixel_column) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                   c   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   b   d       <    else if ((sprite_row + 12 < pixel_row) && (pixel_row < sprite_row  + 15) && ((sprite_column + 3 == pixel_column) || (sprite_column + 3 == pixel_column) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    �   c    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   �   �       ?    else if ((sprite_row + 12 < pixel_row) && (pixel_row < sprite_row  + 15) && ((sprite_column + 22 == pixel_column) || (sprite_column + 23 == pixel_column) || ((sprite_column + 26 < pixel_column) && (pixel_column < sprite_column + 31)) || (pixel_column == sprite_column + 33) || (pixel_column == sprite_column + 34)))5�_�      	              �   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   �   �       ?    else if ((sprite_row + 12 < pixel_row) && (pixel_row < sprite_row  + 15) && ((sprite_column + 23 == pixel_column) || (sprite_column + 23 == pixel_column) || ((sprite_column + 26 < pixel_column) && (pixel_column < sprite_column + 31)) || (pixel_column == sprite_column + 33) || (pixel_column == sprite_column + 34)))5�_�      
           	   �   c    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   �   �       ?    else if ((sprite_row + 12 < pixel_row) && (pixel_row < sprite_row  + 15) && ((sprite_column + 42 == pixel_column) || (sprite_column + 43 == pixel_column) || ((sprite_column + 46 < pixel_column) && (pixel_column < sprite_column + 51)) || (pixel_column == sprite_column + 53) || (pixel_column == sprite_column + 54)))5�_�   	              
   �   �    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   �   �       ?    else if ((sprite_row + 12 < pixel_row) && (pixel_row < sprite_row  + 15) && ((sprite_column + 43 == pixel_column) || (sprite_column + 43 == pixel_column) || ((sprite_column + 46 < pixel_column) && (pixel_column < sprite_column + 51)) || (pixel_column == sprite_column + 53) || (pixel_column == sprite_column + 54)))5�_�   
                 �   �    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   �   �       ?    else if ((sprite_row + 12 < pixel_row) && (pixel_row < sprite_row  + 15) && ((sprite_column + 43 == pixel_column) || (sprite_column + 43 == pixel_column) || ((sprite_column + 46 < pixel_column) && (pixel_column < sprite_column + 51)) || (pixel_column == sprite_column + 53) || (pixel_column == sprite_column + 54)))5�_�                    g       ����                                                                                                                                                                                                                                                                                                                                                             d�(     �   g   i      �   g   h      5�_�                    h       ����                                                                                                                                                                                                                                                                                                                                                             d�+     �   g   i       <    else if ((sprite_row + 12 < pixel_row) && (pixel_row < sprite_row  + 15) && ((sprite_column + 3 == pixel_column) || (sprite_column + 4 == pixel_column) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   J    ����                                                                                                                                                                                                                                                                                                                                                             d�.     �   g   i       <    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 15) && ((sprite_column + 3 == pixel_column) || (sprite_column + 4 == pixel_column) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   `    ����                                                                                                                                                                                                                                                                                                                                                             d�K     �   g   i       <    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 3 == pixel_column) || (sprite_column + 4 == pixel_column) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   `    ����                                                                                                                                                                                                                                                                                                                                                             d�K     �   g   i       ;    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column  3 == pixel_column) || (sprite_column + 4 == pixel_column) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   `    ����                                                                                                                                                                                                                                                                                                                                                             d�K     �   g   i       :    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column 3 == pixel_column) || (sprite_column + 4 == pixel_column) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   _    ����                                                                                                                                                                                                                                                                                                                                                             d�L     �   g   i       9    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column  == pixel_column) || (sprite_column + 4 == pixel_column) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�Q     �   g   i       8    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column == pixel_column) || (sprite_column + 4 == pixel_column) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�Y     �   g   i       8    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column == pixel_column) || (sprite_column + 1 == pixel_column) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   o    ����                                                                                                                                                                                                                                                                                                                                                             d�g     �   g   i       7    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column == pixel_column) || (sprite_column + 1 == pixel_column) || (sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�q     �   g   i       ;    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column == pixel_column + 1) || (sprite_column + 1 == pixel_column) || (sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�r     �   g   i       ;    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column == pixel_column + 1) || (sprite_column +21 == pixel_column) || (sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�s     �   g   i       ;    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column == pixel_column + 1) || (sprite_column +22 == pixel_column) || (sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�t     �   g   i       :    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column == pixel_column + 1) || (sprite_column +2 == pixel_column) || (sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   _    ����                                                                                                                                                                                                                                                                                                                                                             d�{     �   g   i       ;    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column == pixel_column + 1) || (sprite_column + 2 == pixel_column) || (sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   `    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   g   i       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_columni +1 == pixel_column + 1) || (sprite_column + 2 == pixel_column) || (sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   a    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   g   i       >    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column +1 == pixel_column + 1) || (sprite_column + 2 == pixel_column) || (sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   w    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   g   i       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column + 1) || (sprite_column + 2 == pixel_column) || (sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                    h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   g   i       ;    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�                     h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   g   i       <    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 6 x< pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�      !               h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   g   i       <    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 6 == pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�       "           !   h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   g   i       <    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 3 == pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�   !   #           "   h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   g   i       <    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 5 == pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�   "   $           #   h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   g   i       <    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 5 == pixel_column) || (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�   #   %           $   h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   g   i       =    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 5 == pixel_column) || (pixel_column == sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�   $   &           %   h   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   g   i       <    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 5 == pixel_column) || (pixel_column == sprite_column + 6)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�   %   '           &   h      ����                                                                                                                                                                                                                                                                                                                                                             d��     �   g   i       ;    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 5 == pixel_column) || (pixel_column == sprite_column + 6) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5�_�   &   (           '   h  8    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   g   i       ;    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 5 == pixel_column) || (pixel_column == sprite_column + 6) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 14)))5�_�   '   )           (   i       ����                                                                                                                                                                                                                                                                                                                                                             d��     �   h   i             else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && (pixel_column == ((sprite_column + 1) || (sprite_column + 2) || (sprite_column + 5) || (sprite_column + 6) || (sprite_column + 11) || (sprite_column + 12) || (sprite_column + 15) || (sprite_column + 16))))5�_�   (   *           )   �       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   �   �      �   �   �      5�_�   )   +           *   �       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   �   �         !    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && (pixel_column == ((sprite_column + 21) || (sprite_column + 22) || (sprite_column + 25) || (sprite_column + 26) || (sprite_column + 31) || (sprite_column + 32) || (sprite_column + 35) || (sprite_column + 36))))5�_�   *   ,           +   �   b    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   �   �       ;    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 5 == pixel_column) || (pixel_column == sprite_column + 6) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 12)))5�_�   +   -           ,   �   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   �   �       <    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 5 == pixel_column) || (pixel_column == sprite_column + 6) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 12)))5�_�   ,   .           -   �   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   �   �       =    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 5 == pixel_column) || (pixel_column == sprite_column + 6) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 12)))5�_�   -   /           .   �   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   �   �       >    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column +2 5 == pixel_column) || (pixel_column == sprite_column + 6) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 12)))5�_�   .   0           /   �   �    ����                                                                                                                                                                                                                                                                                                                                                             d�      �   �   �       =    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 5 == pixel_column) || (pixel_column == sprite_column + 6) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 12)))5�_�   /   1           0   �   �    ����                                                                                                                                                                                                                                                                                                                                                             d�$     �   �   �       >    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 6) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 12)))5�_�   0   2           1   �      ����                                                                                                                                                                                                                                                                                                                                                             d�&     �   �   �       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 12)))5�_�   1   3           2   �  ;    ����                                                                                                                                                                                                                                                                                                                                                             d�+     �   �   �       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 12)))5�_�   2   4           3   �       ����                                                                                                                                                                                                                                                                                                                                                             d�5     �   �   �      �   �   �      5�_�   3   5           4   �       ����                                                                                                                                                                                                                                                                                                                                                             d�6     �   �   �         !    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && (pixel_column == ((sprite_column + 41) || (sprite_column + 42) || (sprite_column + 45) || (sprite_column + 46) || (sprite_column + 51) || (sprite_column + 52) || (sprite_column + 55) || (sprite_column + 56))))5�_�   4   6           5   �   b    ����                                                                                                                                                                                                                                                                                                                                                             d�<     �   �   �       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 32)))5�_�   5   7           6   �   �    ����                                                                                                                                                                                                                                                                                                                                                             d�?     �   �   �       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 32)))5�_�   6   8           7   �   �    ����                                                                                                                                                                                                                                                                                                                                                             d�A     �   �   �       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 42 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 32)))5�_�   7   9           8   �   �    ����                                                                                                                                                                                                                                                                                                                                                             d�D     �   �   �       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 42 == pixel_column) || (sprite_column + 45 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 32)))5�_�   8   :           9   �      ����                                                                                                                                                                                                                                                                                                                                                             d�F     �   �   �       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 42 == pixel_column) || (sprite_column + 45 == pixel_column) || (pixel_column == sprite_column + 46) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 32)))5�_�   9   ;           :   �      ����                                                                                                                                                                                                                                                                                                                                                             d�H     �   �   �       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 42 == pixel_column) || (sprite_column + 45 == pixel_column) || (pixel_column == sprite_column + 46) || (pixel_column == sprite_column + 41) || (pixel_column == sprite_column + 32)))5�_�   :   <           ;   �  :    ����                                                                                                                                                                                                                                                                                                                                                             d�o     �   �   �       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 42 == pixel_column) || (sprite_column + 45 == pixel_column) || (pixel_column == sprite_column + 46) || (pixel_column == sprite_column + 51) || (pixel_column == sprite_column + 32)))5�_�   ;   =           <   h  9    ����                                                                                                                                                                                                                                                                                                                            h   �       h  8       v  8    d�     �   g   i       ;    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 5 == pixel_column) || (pixel_column == sprite_column + 6) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 12)))5�_�   <   >           =   h  <    ����                                                                                                                                                                                                                                                                                                                            h   �       h  8       v  8    d�     �   g   i       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 5 == pixel_column) || (pixel_column == sprite_column + 6) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 12) || ))�   h   i      5�_�   =   ?           >   h  _    ����                                                                                                                                                                                                                                                                                                                            h   �       h  8       v  8    d�     �   g   i       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 5 == pixel_column) || (pixel_column == sprite_column + 6) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 12) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 12)))5�_�   >   @           ?   h  �    ����                                                                                                                                                                                                                                                                                                                            h   �       h  8       v  8    d�     �   g   i       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 1 == pixel_column) || (sprite_column + 2 == pixel_column) || (sprite_column + 5 == pixel_column) || (pixel_column == sprite_column + 6) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 12) || (pixel_column == sprite_column + 15) || (pixel_column == sprite_column + 12)))5�_�   ?   A           @   �  =    ����                                                                                                                                                                                                                                                                                                                            h  :       h  �       v  �    d��     �   �   �       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 32)))�   �   �      5�_�   @   B           A   �  =    ����                                                                                                                                                                                                                                                                                                                            h  :       h  �       v  �    d��     �   �   �       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 32))|| (pixel_column == sprite_column + 15) || (pixel_column == sprite_column + 16))5�_�   A   C           B   �  =    ����                                                                                                                                                                                                                                                                                                                            h  :       h  �       v  �    d��     �   �   �       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 32)|| (pixel_column == sprite_column + 15) || (pixel_column == sprite_column + 16))5�_�   B   D           C   �  b    ����                                                                                                                                                                                                                                                                                                                            h  :       h  �       v  �    d��     �   �   �       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 32) || (pixel_column == sprite_column + 15) || (pixel_column == sprite_column + 16))5�_�   C   E           D   �  d    ����                                                                                                                                                                                                                                                                                                                            h  :       h  �       v  �    d��     �   �   �       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 32) || (pixel_column == sprite_column + r315) || (pixel_column == sprite_column + 16))5�_�   D   F           E   �  c    ����                                                                                                                                                                                                                                                                                                                            h  :       h  �       v  �    d��     �   �   �       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 32) || (pixel_column == sprite_column + 15) || (pixel_column == sprite_column + 16))5�_�   E   G           F   �  �    ����                                                                                                                                                                                                                                                                                                                            h  :       h  �       v  �    d��     �   �   �       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 32) || (pixel_column == sprite_column + 35) || (pixel_column == sprite_column + 16))5�_�   F   J           G   �  �    ����                                                                                                                                                                                                                                                                                                                            h  :       h  �       v  �    d��     �   �   �       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 21 == pixel_column) || (sprite_column + 22 == pixel_column) || (sprite_column + 25 == pixel_column) || (pixel_column == sprite_column + 26) || (pixel_column == sprite_column + 31) || (pixel_column == sprite_column + 32) || (pixel_column == sprite_column + 35) || (pixel_column == sprite_column + 36))5�_�   G   K   I       J   �  <    ����                                                                                                                                                                                                                                                                                                                            �  <       �   �       v   �    d�G     �   �   �       ?    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 42 == pixel_column) || (sprite_column + 45 == pixel_column) || (pixel_column == sprite_column + 46) || (pixel_column == sprite_column + 51) || (pixel_column == sprite_column + 52)))�   �   �      5�_�   J   L           K   �  =    ����                                                                                                                                                                                                                                                                                                                            �  <       �   �       v   �    d�O     �   �   �       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 42 == pixel_column) || (sprite_column + 45 == pixel_column) || (pixel_column == sprite_column + 46) || (pixel_column == sprite_column + 51) || (pixel_column == sprite_column + 52)|| (pixel_column == sprite_column + 51) || (pixel_column == sprite_column + 52)))5�_�   K   M           L   �  c    ����                                                                                                                                                                                                                                                                                                                            �  <       �   �       v   �    d�W     �   �   �       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 42 == pixel_column) || (sprite_column + 45 == pixel_column) || (pixel_column == sprite_column + 46) || (pixel_column == sprite_column + 51) || (pixel_column == sprite_column + 52) || (pixel_column == sprite_column + 51) || (pixel_column == sprite_column + 52)))5�_�   L   N           M   �  e    ����                                                                                                                                                                                                                                                                                                                            �  <       �   �       v   �    d�X     �   �   �       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 42 == pixel_column) || (sprite_column + 45 == pixel_column) || (pixel_column == sprite_column + 46) || (pixel_column == sprite_column + 51) || (pixel_column == sprite_column + 52) || (pixel_column == sprite_column + 551) || (pixel_column == sprite_column + 52)))5�_�   M               N   �  �    ����                                                                                                                                                                                                                                                                                                                            �  <       �   �       v   �    d�\    �   �   �       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 42 == pixel_column) || (sprite_column + 45 == pixel_column) || (pixel_column == sprite_column + 46) || (pixel_column == sprite_column + 51) || (pixel_column == sprite_column + 52) || (pixel_column == sprite_column + 55) || (pixel_column == sprite_column + 52)))5�_�   G       H   J   I   �  =    ����                                                                                                                                                                                                                                                                                                                            �  <       �   �       v   �    d�C     �   �   �      �   �   �       �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 42 == pixel_column) || (sprite_column + 45 == pixel_column) || (pixel_column == sprite_column + 46) || (pixel_column == sprite_column + 51) || (pixel_column == sprite_column + 52))|| (pixel_column == sprite_column + 51) || (pixel_column == sprite_column + 52))5�_�   G           I   H   �  =    ����                                                                                                                                                                                                                                                                                                                            h  :       h  �       v  �    d�)     �   �   �      �   �   �       @    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && ((sprite_column + 41 == pixel_column) || (sprite_column + 42 == pixel_column) || (sprite_column + 45 == pixel_column) || (pixel_column == sprite_column + 46) || (pixel_column == sprite_column + 51) || (pixel_column == sprite_column + 52))))5�_�                    c   �    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   b   d       <    else if ((sprite_row + 12 < pixel_row) && (pixel_row < sprite_row  + 15) && ((sprite_column + 3 == pixel_column) || (sprite_column + 4 == pixel_column) || ((sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11)) || (pixel_column == sprite_column + 13) || (pixel_column == sprite_column + 14)))5��