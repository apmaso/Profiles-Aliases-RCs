Vim�UnDo� �j�~1���L��!���u�Չ�M[��fRͪ�   A                                   dw    _�                             ����                                                                                                                                                                                                                                                                                                                                                             dk     �                "    output wire  [11:0] btn_row_o,5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             dq     �                logic [11:0] btn_row_reg;5�_�                              ����                                                                                                                                                                                                                                                                                                                                                             dv    �                 btn_row_reg = 460;5��