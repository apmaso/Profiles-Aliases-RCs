Vim�UnDo� b�v�83���^>B��=�1��C�#9C�$   �  �	else if ((sprite_row + 230 < pixel_row) && (pixel_row < sprite_row + 241) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))   q                      d�    _�                    9        ����                                                                                                                                                                                                                                                                                                                                                             d
     �   8   D   �      	// Row 51 - 100�   9   :   �    5�_�                    9        ����                                                                                                                                                                                                                                                                                                                                                             d     �   8   :   �      		// Row 51 - 905�_�                    C        ����                                                                                                                                                                                                                                                                                                                                                             dC     �   B   C          // Row 51 - 1005�_�                    C       ����                                                                                                                                                                                                                                                                                                                                                             dD     �   B   C         �    else if ((sprite_row + 50 < pixel_row) && (pixel_row < sprite_row + 101) && (((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 210 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    C       ����                                                                                                                                                                                                                                                                                                                                                             dD     �   B   C                  begin5�_�      	              C       ����                                                                                                                                                                                                                                                                                                                                                             dE     �   B   C                       loser_pix = 4'b1111;5�_�      
           	   C       ����                                                                                                                                                                                                                                                                                                                                                             dE     �   B   C                  end5�_�   	              
   D   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 91)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   
                 D   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 0 < pixel_column) && (pixel_column < sprite_column + 91)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 91)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + xi1391)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + xi131)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D   �    ����                                                                                                                                                                                                                                                                                                                                                             d	     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D   �    ����                                                                                                                                                                                                                                                                                                                                                             d     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  6    ����                                                                                                                                                                                                                                                                                                                                                             d     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  4    ����                                                                                                                                                                                                                                                                                                                                                             d     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  Q    ����                                                                                                                                                                                                                                                                                                                                                             d     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  �    ����                                                                                                                                                                                                                                                                                                                                                             d'     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  �    ����                                                                                                                                                                                                                                                                                                                                                             d/     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  �    ����                                                                                                                                                                                                                                                                                                                                                             d/     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))|| ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  �    ����                                                                                                                                                                                                                                                                                                                                                             d/     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))| ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  �    ����                                                                                                                                                                                                                                                                                                                                                             d/     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  �    ����                                                                                                                                                                                                                                                                                                                                                             d/     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  �    ����                                                                                                                                                                                                                                                                                                                                                             d/     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))(sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))prite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))rite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))ite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                     D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))te_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�      !               D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))e_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�       "           !   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   !   #           "   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   "   $           #   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))olumn + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   #   %           $   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))lumn + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   $   &           %   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))umn + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   %   '           &   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))mn + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   &   (           '   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))n + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   '   )           (   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   (   *           )   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))+ 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   )   +           *   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   *   ,           +   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   +   -           ,   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))70 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   ,   .           -   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))0 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   -   /           .   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   .   0           /   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))< pixel_column) && (pixel_column < sprite_column + 281))))5�_�   /   1           0   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) pixel_column) && (pixel_column < sprite_column + 281))))5�_�   0   2           1   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))pixel_column) && (pixel_column < sprite_column + 281))))5�_�   1   3           2   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))ixel_column) && (pixel_column < sprite_column + 281))))5�_�   2   4           3   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))xel_column) && (pixel_column < sprite_column + 281))))5�_�   3   5           4   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))el_column) && (pixel_column < sprite_column + 281))))5�_�   4   6           5   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))l_column) && (pixel_column < sprite_column + 281))))5�_�   5   7           6   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))_column) && (pixel_column < sprite_column + 281))))5�_�   6   8           7   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))column) && (pixel_column < sprite_column + 281))))5�_�   7   9           8   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))olumn) && (pixel_column < sprite_column + 281))))5�_�   8   :           9   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))lumn) && (pixel_column < sprite_column + 281))))5�_�   9   ;           :   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))umn) && (pixel_column < sprite_column + 281))))5�_�   :   <           ;   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d0     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))mn) && (pixel_column < sprite_column + 281))))5�_�   ;   =           <   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d1     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))n) && (pixel_column < sprite_column + 281))))5�_�   <   >           =   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d1     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))) && (pixel_column < sprite_column + 281))))5�_�   =   ?           >   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d1     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) && (pixel_column < sprite_column + 281))))5�_�   >   @           ?   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d1     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))&& (pixel_column < sprite_column + 281))))5�_�   ?   A           @   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d1     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))& (pixel_column < sprite_column + 281))))5�_�   @   B           A   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d1     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) (pixel_column < sprite_column + 281))))5�_�   A   C           B   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d1     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))(pixel_column < sprite_column + 281))))5�_�   B   D           C   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d1     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))pixel_column < sprite_column + 281))))5�_�   C   E           D   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d1     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))ixel_column < sprite_column + 281))))5�_�   D   F           E   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d1     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))xel_column < sprite_column + 281))))5�_�   E   G           F   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d1     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))el_column < sprite_column + 281))))5�_�   F   H           G   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d1     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))l_column < sprite_column + 281))))5�_�   G   I           H   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))_column < sprite_column + 281))))5�_�   H   J           I   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))column < sprite_column + 281))))5�_�   I   K           J   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))olumn < sprite_column + 281))))5�_�   J   L           K   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))lumn < sprite_column + 281))))5�_�   K   M           L   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))umn < sprite_column + 281))))5�_�   L   N           M   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))mn < sprite_column + 281))))5�_�   M   O           N   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))n < sprite_column + 281))))5�_�   N   P           O   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) < sprite_column + 281))))5�_�   O   Q           P   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))< sprite_column + 281))))5�_�   P   R           Q   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) sprite_column + 281))))5�_�   Q   S           R   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))sprite_column + 281))))5�_�   R   T           S   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))prite_column + 281))))5�_�   S   U           T   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))rite_column + 281))))5�_�   T   V           U   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))ite_column + 281))))5�_�   U   W           V   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))te_column + 281))))5�_�   V   X           W   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))e_column + 281))))5�_�   W   Y           X   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))_column + 281))))5�_�   X   Z           Y   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))column + 281))))5�_�   Y   [           Z   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))olumn + 281))))5�_�   Z   \           [   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))lumn + 281))))5�_�   [   ]           \   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d2     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))umn + 281))))5�_�   \   ^           ]   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d3     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))mn + 281))))5�_�   ]   _           ^   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d3     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))n + 281))))5�_�   ^   `           _   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d3     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) + 281))))5�_�   _   a           `   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d3     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))+ 281))))5�_�   `   b           a   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d3     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) 281))))5�_�   a   c           b   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d3     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))281))))5�_�   b   d           c   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d4     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))81))))5�_�   c   e           d   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d4     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))1))))5�_�   d   f           e   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d4     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))))))5�_�   e   g           f   D  �    ����                                                                                                                                                                                                                                                                                                                                                             d5     �   C   E   �     �	else if ((sprite_row + 150 < pixel_row) && (pixel_row < sprite_row + 161) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)))))5�_�   f   h           g   H       ����                                                                                                                                                                                                                                                                                                                                                             dv     �   G   I   �      	// Rows 161 - 1805�_�   g   i           h   I   G    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     1	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 181) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 91)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 220 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   h   l           i   I   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     1	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 91)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 220 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   i   m   j       l   I   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     1	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 91)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 220 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   l   n           m   I   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     1	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 220 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   m   o           n   I  4    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     1	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 220 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   n   p           o   I  N    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     1	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 220 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   o   q           p   I  N    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     0	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 00 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 220 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   p   r           q   I  N    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     /	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 0 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 220 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   q   s           r   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     1	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 220 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   r   t           s   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     1	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 220 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   s   u           t   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     2	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 2320 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   t   v           u   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     1	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   u   w           v   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     1	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   v   x           w   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     0	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))|| ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   w   y           x   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     /	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))| ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   x   z           y   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     .	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   y   {           z   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     -	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   z   |           {   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     ,	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))(sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   {   }           |   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     +	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   |   ~           }   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     *	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))prite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   }              ~   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     )	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))rite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   ~   �              I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     (	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))ite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�      �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     '	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))te_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     &	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))e_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     %	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     $	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     #	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))olumn + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     "	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))lumn + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     !	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))umn + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �      	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))mn + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))n + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))+ 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))70 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))0 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))< pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))ixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))xel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))el_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))l_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))olumn) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))lumn) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))umn) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))mn) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     
	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))n) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     		else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))&& (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))& (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) (pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))(pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))pixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))ixel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))xel_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �      	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))el_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))l_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))_column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))column < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))olumn < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))lumn < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))umn < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))mn < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))n < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) < sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))< sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))sprite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))prite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))rite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))ite_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))te_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))e_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))_column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))column + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))olumn + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))lumn + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))umn + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))mn + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))n + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) + 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))+ 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)) 281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))281))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))81))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))1))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281)))))5�_�   �   �           �   I  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   M   	    ����                                                                                                                                                                                                                                                                                                                                                             d     �   L   N   �      	// Rows 181 - 2005�_�   �   �           �   M   	    ����                                                                                                                                                                                                                                                                                                                                                             d     �   L   N   �      	// Rows 81 - 2005�_�   �   �           �   M   	    ����                                                                                                                                                                                                                                                                                                                                                             d     �   L   N   �      	// Rows 1 - 2005�_�   �   �           �   M   	    ����                                                                                                                                                                                                                                                                                                                                                             d     �   L   N   �      	// Rows  - 2005�_�   �   �           �   M   	    ����                                                                                                                                                                                                                                                                                                                                                             d     �   L   N   �      	// Rows - 2005�_�   �   �           �   M   	    ����                                                                                                                                                                                                                                                                                                                                                             d     �   L   N   �      	// Rows  2005�_�   �   �           �   M   	    ����                                                                                                                                                                                                                                                                                                                                                             d     �   L   N   �      	// Rows 2005�_�   �   �           �   M   	    ����                                                                                                                                                                                                                                                                                                                                                             d     �   L   N   �      	// Rows 005�_�   �   �           �   M   	    ����                                                                                                                                                                                                                                                                                                                                                             d     �   L   N   �      
	// Rows 05�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                                                             d     �   L   N   �      		// Rows 5�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                                                             d     �   L   N   �      	// Rows�   M   N   �    5�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                                                             d     �   M   O   �    �   M   N   �    5�_�   �   �           �   O       ����                                                                                                                                                                                                                                                                                                                                                             d     �   N   O         6	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 201) && (((sprite_column + 10 < pixel_column) && (pixel_column < sprite_column + 21)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                                                             d      �   L   N   �      		// Rows 5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                                                             d(     �   M   O   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�   �   �           �   N   H    ����                                                                                                                                                                                                                                                                                                                                                             d/     �   M   O   �     �	else if ((sprite_row + 170 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�   �   �           �   N  4    ����                                                                                                                                                                                                                                                                                                                                                             dU     �   M   O   �     �	else if ((sprite_row + 170 < pixel_row) && (pixel_row < sprite_row + 181) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�   �   �           �   N  7    ����                                                                                                                                                                                                                                                                                                                                                             dW     �   M   O   �     �	else if ((sprite_row + 170 < pixel_row) && (pixel_row < sprite_row + 181) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 1r321)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�   �   �           �   I  5    ����                                                                                                                                                                                                                                                                                                                                                             dY     �   H   J   �     �	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�   �   �           �   N  P    ����                                                                                                                                                                                                                                                                                                                                                             d}     �   M   O   �     �	else if ((sprite_row + 170 < pixel_row) && (pixel_row < sprite_row + 181) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�   �   �           �   N  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   M   O   �     �	else if ((sprite_row + 170 < pixel_row) && (pixel_row < sprite_row + 181) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 161)) ||  ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   Q   S   �      	// Rows 201 - 2105�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   Q   S   �      	// Rows201 - 2105�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   Q   S   �      	// Rows01 - 2105�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   Q   S   �      	// Rows1 - 2105�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   Q   S   �      	// Rows - 2105�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   Q   S   �      	// Rows- 2105�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   Q   S   �      	// Rows 2105�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   Q   S   �      	// Rows2105�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   Q   S   �      
	// Rows105�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   Q   S   �      		// Rows05�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   Q   S   �      	// Rows5�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   Q   S   �      	// Rows5�_�   �   �           �   S       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   R   T   �     5	else if ((sprite_row + 200 < pixel_row) && (pixel_row < sprite_row + 211) && (((sprite_column + 10 < pixel_column) && (pixel_column < sprite_column + 21)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S   I    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   R   T   �     5	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 211) && (((sprite_column + 10 < pixel_column) && (pixel_column < sprite_column + 21)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S   I    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   R   T   �     5	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 195) && (((sprite_column + 10 < pixel_column) && (pixel_column < sprite_column + 21)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S   c    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   R   T   �     5	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column + 10 < pixel_column) && (pixel_column < sprite_column + 21)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   R   T   �     0	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 21)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   R   T   �     0	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  5    ����                                                                                                                                                                                                                                                                                                                                                             d     �   R   T   �     0	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  Q    ����                                                                                                                                                                                                                                                                                                                                                             d     �   R   T   �     0	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             d     �   R   T   �     0	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             d@     �   R   T   �     0	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dH     �   R   T   �     0	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dK     �   R   T   �     0	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     0	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     /	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))|| ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     .	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))| ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     -	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     ,	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     +	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))(sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     *	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     )	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))prite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �   �           �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     (	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))rite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �              �   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     '	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))ite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   �                S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     &	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))te_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                  S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     %	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))e_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     $	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     #	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dN     �   R   T   �     "	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))olumn + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     !	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))lumn + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �      	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))umn + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))mn + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�    	             S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))n + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�    
          	   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  	            
   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))+ 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  
               S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))70 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))0 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))< pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))pixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))ixel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))xel_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))el_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))l_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))_column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))column) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))olumn) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))lumn) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))umn) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     
	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))mn) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     		else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))n) && (pixel_column < sprite_column + 281))))5�_�                 S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))) && (pixel_column < sprite_column + 281))))5�_�                  S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) && (pixel_column < sprite_column + 281))))5�_�    !              S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))&& (pixel_column < sprite_column + 281))))5�_�     "          !   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))& (pixel_column < sprite_column + 281))))5�_�  !  #          "   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) (pixel_column < sprite_column + 281))))5�_�  "  $          #   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))(pixel_column < sprite_column + 281))))5�_�  #  %          $   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))pixel_column < sprite_column + 281))))5�_�  $  &          %   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �     	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))ixel_column < sprite_column + 281))))5�_�  %  '          &   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dO     �   R   T   �      	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))xel_column < sprite_column + 281))))5�_�  &  (          '   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))el_column < sprite_column + 281))))5�_�  '  )          (   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))l_column < sprite_column + 281))))5�_�  (  *          )   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))_column < sprite_column + 281))))5�_�  )  +          *   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))column < sprite_column + 281))))5�_�  *  ,          +   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))olumn < sprite_column + 281))))5�_�  +  -          ,   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))lumn < sprite_column + 281))))5�_�  ,  .          -   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))umn < sprite_column + 281))))5�_�  -  /          .   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))mn < sprite_column + 281))))5�_�  .  0          /   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))n < sprite_column + 281))))5�_�  /  1          0   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) < sprite_column + 281))))5�_�  0  2          1   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))< sprite_column + 281))))5�_�  1  3          2   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) sprite_column + 281))))5�_�  2  4          3   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))sprite_column + 281))))5�_�  3  5          4   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))prite_column + 281))))5�_�  4  6          5   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))rite_column + 281))))5�_�  5  7          6   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))ite_column + 281))))5�_�  6  8          7   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))te_column + 281))))5�_�  7  9          8   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))e_column + 281))))5�_�  8  :          9   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))_column + 281))))5�_�  9  ;          :   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))column + 281))))5�_�  :  <          ;   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))olumn + 281))))5�_�  ;  =          <   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))lumn + 281))))5�_�  <  >          =   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))umn + 281))))5�_�  =  ?          >   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))mn + 281))))5�_�  >  @          ?   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))n + 281))))5�_�  ?  A          @   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dP     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) + 281))))5�_�  @  B          A   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dQ     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))+ 281))))5�_�  A  C          B   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dQ     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)) 281))))5�_�  B  D          C   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dQ     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))281))))5�_�  C  E          D   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dQ     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))81))))5�_�  D  F          E   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dR     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))1))))5�_�  E  G          F   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dR     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))))5�_�  F  H          G   S  �    ����                                                                                                                                                                                                                                                                                                                                                             dR     �   R   T   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241)))))5�_�  G  I          H   W   	    ����                                                                                                                                                                                                                                                                                                                                                             da     �   V   X   �      	// Rows 211 - 2205�_�  H  J          I   W   	    ����                                                                                                                                                                                                                                                                                                                                                             da     �   V   X   �      	// Rows 11 - 2205�_�  I  K          J   W   	    ����                                                                                                                                                                                                                                                                                                                                                             da     �   V   X   �      	// Rows 1 - 2205�_�  J  L          K   W   	    ����                                                                                                                                                                                                                                                                                                                                                             da     �   V   X   �      	// Rows  - 2205�_�  K  M          L   W   	    ����                                                                                                                                                                                                                                                                                                                                                             db     �   V   X   �      	// Rows - 2205�_�  L  N          M   W   	    ����                                                                                                                                                                                                                                                                                                                                                             db     �   V   X   �      	// Rows  2205�_�  M  O          N   W   	    ����                                                                                                                                                                                                                                                                                                                                                             db     �   V   X   �      	// Rows 2205�_�  N  P          O   W   	    ����                                                                                                                                                                                                                                                                                                                                                             db     �   V   X   �      	// Rows 205�_�  O  Q          P   W   	    ����                                                                                                                                                                                                                                                                                                                                                             db     �   V   X   �      
	// Rows 05�_�  P  R          Q   W       ����                                                                                                                                                                                                                                                                                                                                                             d}     �   V   X   �      		// Rows 5�_�  Q  S          R   X       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   W   Y   �     �	else if ((sprite_row + 210 < pixel_row) && (pixel_row < sprite_row + 221) && (((sprite_column + 20 < pixel_column) && (pixel_column < sprite_column + 31)) || ((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 60 < pixel_column) && (pixel_column < sprite_column + 71)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  R  T          S   X       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   W   Y   �     �	else if ((sprite_row + xx210 < pixel_row) && (pixel_row < sprite_row + 221) && (((sprite_column + 20 < pixel_column) && (pixel_column < sprite_column + 31)) || ((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 60 < pixel_column) && (pixel_column < sprite_column + 71)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  S  U          T   X       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   W   Y   �     �	else if ((sprite_row + 196 < pixel_row) && (pixel_row < sprite_row + 221) && (((sprite_column + 20 < pixel_column) && (pixel_column < sprite_column + 31)) || ((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 60 < pixel_column) && (pixel_column < sprite_column + 71)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  T  V          U   X   H    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   W   Y   �     �	else if ((sprite_row + 195 < pixel_row) && (pixel_row < sprite_row + 221) && (((sprite_column + 20 < pixel_column) && (pixel_column < sprite_column + 31)) || ((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 60 < pixel_column) && (pixel_column < sprite_column + 71)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  U  W          V   W       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   W   Y   �    �   W   X   �    5�_�  V  X          W   Y       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   X   Y         �	else if ((sprite_row + 195 < pixel_row) && (pixel_row < sprite_row + 201) && (((sprite_column + 20 < pixel_column) && (pixel_column < sprite_column + 31)) || ((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 60 < pixel_column) && (pixel_column < sprite_column + 71)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  W  Y          X   X       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   W   Y   �     �	else if ((sprite_row + 180 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  X  Z          Y   X       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   W   Y   �     �	else if ((sprite_row + 190 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  Y  \          Z   X   I    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   W   Y   �     �	else if ((sprite_row + 195 < pixel_row) && (pixel_row < sprite_row + 196) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  Z  ]  [      \   X  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   W   Y   �     �	else if ((sprite_row + 195 < pixel_row) && (pixel_row < sprite_row + 201) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  \  ^          ]   \   	    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   [   ]   �      	// Rows 221 - 2305�_�  ]  _          ^   \   	    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   [   ]   �      	// Rows 21 - 2305�_�  ^  `          _   \   	    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   [   ]   �      	// Rows 1 - 2305�_�  _  a          `   \   	    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   [   ]   �      	// Rows  - 2305�_�  `  b          a   \   	    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   [   ]   �      	// Rows - 2305�_�  a  c          b   \   	    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   [   ]   �      	// Rows  2305�_�  b  d          c   \   	    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   [   ]   �      	// Rows 2305�_�  c  e          d   \   	    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   [   ]   �      	// Rows 305�_�  d  f          e   \   	    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   [   ]   �      
	// Rows 05�_�  e  g          f   \       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   [   ]   �      	// Rows 205�_�  f  h          g   ]       ����                                                                                                                                                                                                                                                                                                                                                             d     �   \   ]         �	else if ((sprite_row + 220 < pixel_row) && (pixel_row < sprite_row + 231) && (((sprite_column + 20 < pixel_column) && (pixel_column < sprite_column + 31)) || ((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 60 < pixel_column) && (pixel_column < sprite_column + 71)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 250 < pixel_column) && (pixel_column < sprite_column + 261)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  g  i          h   \       ����                                                                                                                                                                                                                                                                                                                                                             d	     �   \   ^   �    �   \   ]   �    5�_�  h  j          i   \       ����                                                                                                                                                                                                                                                                                                                                                             d     �   \   ^   �    �   \   ]   �    5�_�  i  k          j   ^       ����                                                                                                                                                                                                                                                                                                                                                             d     �   ]   ^         �	else if ((sprite_row + 220 < pixel_row) && (pixel_row < sprite_row + 231) && (((sprite_column + 20 < pixel_column) && (pixel_column < sprite_column + 31)) || ((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 60 < pixel_column) && (pixel_column < sprite_column + 71)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 250 < pixel_column) && (pixel_column < sprite_column + 261)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  j  l          k   ]       ����                                                                                                                                                                                                                                                                                                                                                             d     �   \   ^   �     �	else if ((sprite_row + 195 < pixel_row) && (pixel_row < sprite_row + 201) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 261))))5�_�  k  m          l   ]   I    ����                                                                                                                                                                                                                                                                                                                                                             d!     �   \   ^   �     �	else if ((sprite_row + 200 < pixel_row) && (pixel_row < sprite_row + 201) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 261))))5�_�  l  n          m   ]  O    ����                                                                                                                                                                                                                                                                                                                                                             d;     �   \   ^   �     �	else if ((sprite_row + 200 < pixel_row) && (pixel_row < sprite_row + 206) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 261))))5�_�  m  o          n   ]  Q    ����                                                                                                                                                                                                                                                                                                                                                             d=     �   \   ^   �     �	else if ((sprite_row + 200 < pixel_row) && (pixel_row < sprite_row + 206) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 1r70 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 261))))5�_�  n  p          o   ]  �    ����                                                                                                                                                                                                                                                                                                                                                             dB     �   \   ^   �     �	else if ((sprite_row + 200 < pixel_row) && (pixel_row < sprite_row + 206) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 180 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 261))))5�_�  o  q          p   b       ����                                                                                                                                                                                                                                                                                                                                                             d_     �   a   c   �     6	else if ((sprite_row + 230 < pixel_row) && (pixel_row < sprite_row + 241) && (((sprite_column + 30 < pixel_column) && (pixel_column < sprite_column + 41)) || ((sprite_column + 50 < pixel_column) && (pixel_column < sprite_column + 61)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 250 < pixel_column) && (pixel_column < sprite_column + 261)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  p  r          q   a       ����                                                                                                                                                                                                                                                                                                                                                             de     �   `   b   �      	// Rows 231 - 2405�_�  q  s          r   b   H    ����                                                                                                                                                                                                                                                                                                                                                             dn     �   a   c   �     6	else if ((sprite_row + 205 < pixel_row) && (pixel_row < sprite_row + 241) && (((sprite_column + 30 < pixel_column) && (pixel_column < sprite_column + 41)) || ((sprite_column + 50 < pixel_column) && (pixel_column < sprite_column + 61)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 250 < pixel_column) && (pixel_column < sprite_column + 261)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  r  t          s   a       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   a   c   �    �   a   b   �    5�_�  s  u          t   c       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   b   c         6	else if ((sprite_row + 205 < pixel_row) && (pixel_row < sprite_row + 221) && (((sprite_column + 30 < pixel_column) && (pixel_column < sprite_column + 41)) || ((sprite_column + 50 < pixel_column) && (pixel_column < sprite_column + 61)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 250 < pixel_column) && (pixel_column < sprite_column + 261)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  t  v          u   b       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   a   c   �     �	else if ((sprite_row + 200 < pixel_row) && (pixel_row < sprite_row + 206) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 180 < pixel_column) && (pixel_column < sprite_column + 191)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 261))))5�_�  u  w          v   b   G    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   a   c   �     �	else if ((sprite_row + 205 < pixel_row) && (pixel_row < sprite_row + 206) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 180 < pixel_column) && (pixel_column < sprite_column + 191)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 261))))5�_�  v  x          w   b   H    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   a   c   �     �	else if ((sprite_row + 205 < pixel_row) && (pixel_row < sprite_row + 226) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 180 < pixel_column) && (pixel_column < sprite_column + 191)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 261))))5�_�  w  y          x   b  �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   a   c   �     �	else if ((sprite_row + 205 < pixel_row) && (pixel_row < sprite_row + 221) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 180 < pixel_column) && (pixel_column < sprite_column + 191)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 261))))5�_�  x  z          y   f       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   f   h   �    �   f   g   �    5�_�  y  {          z   f   
    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   e   g   �      	// Rows 241 - 2505�_�  z  |          {   f       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   e   g   �      	// Rows 221 - 2505�_�  {  }          |   h       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   g   h         �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column + 30 < pixel_column) && (pixel_column < sprite_column + 41)) || ((sprite_column + 50 < pixel_column) && (pixel_column < sprite_column + 61)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 260 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  |  ~          }   g       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   f   h   �     �	else if ((sprite_row + 205 < pixel_row) && (pixel_row < sprite_row + 221) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 180 < pixel_column) && (pixel_column < sprite_column + 191)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  }            ~   g       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   f   h   �     �	else if ((sprite_row + 225 < pixel_row) && (pixel_row < sprite_row + 221) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 180 < pixel_column) && (pixel_column < sprite_column + 191)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  ~  �             g       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   f   h   �     �	else if ((sprite_row + 221 < pixel_row) && (pixel_row < sprite_row + 221) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 180 < pixel_column) && (pixel_column < sprite_column + 191)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�    �          �   g   G    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   f   h   �     �	else if ((sprite_row + 220 < pixel_row) && (pixel_row < sprite_row + 221) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 180 < pixel_column) && (pixel_column < sprite_column + 191)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   g  O    ����                                                                                                                                                                                                                                                                                                                                                             d	     �   f   h   �     �	else if ((sprite_row + 220 < pixel_row) && (pixel_row < sprite_row + 231) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 180 < pixel_column) && (pixel_column < sprite_column + 191)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   g  �    ����                                                                                                                                                                                                                                                                                                                                                             d     �   f   h   �     �	else if ((sprite_row + 220 < pixel_row) && (pixel_row < sprite_row + 231) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 190 < pixel_column) && (pixel_column < sprite_column + 191)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   g  �    ����                                                                                                                                                                                                                                                                                                                                                             d     �   f   h   �     �	else if ((sprite_row + 220 < pixel_row) && (pixel_row < sprite_row + 231) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 190 < pixel_column) && (pixel_column < sprite_column + 91)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   g  �    ����                                                                                                                                                                                                                                                                                                                                                             d     �   f   h   �     �	else if ((sprite_row + 220 < pixel_row) && (pixel_row < sprite_row + 231) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 190 < pixel_column) && (pixel_column < sprite_column + 1)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   j       ����                                                                                                                                                                                                                                                                                                                            j          e          v  �    d'     �   i   p   �      		end�   j   k   �    5�_�  �  �          �   k   
    ����                                                                                                                                                                                                                                                                                                                            j          e          v  �    d+     �   j   l   �      	// Rows 221 - 2305�_�  �  �          �   k       ����                                                                                                                                                                                                                                                                                                                            j          e          v  �    d.     �   j   l   �      	// Rows 231 - 2305�_�  �  �          �   l       ����                                                                                                                                                                                                                                                                                                                            j          e          v  �    d0     �   k   m   �     �	else if ((sprite_row + 220 < pixel_row) && (pixel_row < sprite_row + 231) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 190 < pixel_column) && (pixel_column < sprite_column + 201)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   l   G    ����                                                                                                                                                                                                                                                                                                                            j          e          v  �    d4     �   k   m   �     �	else if ((sprite_row + 230 < pixel_row) && (pixel_row < sprite_row + 231) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 190 < pixel_column) && (pixel_column < sprite_column + 201)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   l  N    ����                                                                                                                                                                                                                                                                                                                            j          e          v  �    dQ     �   k   m   �     �	else if ((sprite_row + 230 < pixel_row) && (pixel_row < sprite_row + 241) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 190 < pixel_column) && (pixel_column < sprite_column + 201)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   l  N    ����                                                                                                                                                                                                                                                                                                                            j          e          v  �    dQ     �   k   m   �     �	else if ((sprite_row + 230 < pixel_row) && (pixel_row < sprite_row + 241) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 90 < pixel_column) && (pixel_column < sprite_column + 201)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   l  N    ����                                                                                                                                                                                                                                                                                                                            j          e          v  �    dS     �   k   m   �     �	else if ((sprite_row + 230 < pixel_row) && (pixel_row < sprite_row + 241) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 0 < pixel_column) && (pixel_column < sprite_column + 201)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   l  �    ����                                                                                                                                                                                                                                                                                                                            j          e          v  �    dW     �   k   m   �     �	else if ((sprite_row + 230 < pixel_row) && (pixel_row < sprite_row + 241) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 201)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   p        ����                                                                                                                                                                                                                                                                                                                            k           o          v       dw     �   o   v   �      	else�   p   q   �    5�_�  �  �          �   p       ����                                                                                                                                                                                                                                                                                                                            k           o          v       d{     �   o   q   �      		// Rows 231 - 2405�_�  �  �          �   p       ����                                                                                                                                                                                                                                                                                                                            k           o          v       d     �   o   q   �          // Rows 231 - 2405�_�  �  �          �   p       ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   o   q   �          // Rows 241 - 2405�_�  �  �          �   q       ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 230 < pixel_row) && (pixel_row < sprite_row + 241) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   H    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 241) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �  �      �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&(pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&ixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&xel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&el_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&l_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&olumn < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&lumn < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&umn < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&mn < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&n < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&< sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&prite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&rite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&ite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&te_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&e_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&olumn + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&lumn + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&umn + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&mn + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&n + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&+ 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&1)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&|| ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&| ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&(sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&prite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&rite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&ite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&te_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&e_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&olumn + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&lumn + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&umn + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&mn + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&n + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&+ 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&20 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&0 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �             �   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&< pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �                q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                  q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&ixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&xel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&el_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&l_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�    	             q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&olumn) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�    
          	   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&lumn) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  	            
   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&umn) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  
               q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&mn) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&n) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&&& (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&& (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�               q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 00 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 0 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column +  < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                   q  �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�    �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 150 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�               q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&(pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                 q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�                   q   �    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 70 < pixel_column) &&ixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �      �  �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && `(pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && ixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && xel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && el_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && l_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && _column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && olumn < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && lumn < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && umn < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && mn < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && n < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) &&  < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) &&  sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && prite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && rite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && ite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && te_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && e_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && _column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && olumn + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && lumn + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && umn + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && mn + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && n + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) &&  + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) &&  11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && 1)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && )) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && ) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) &&  || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && | ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) &&  ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �  �          �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  �              �   q   r    ����                                                                                                                                                                                                                                                                                                                            k           o          v       d�     �   p   r   �     �	else if ((sprite_row + 240 < pixel_row) && (pixel_row < sprite_row + 251) && (((sprite_column < pixel_column) && (sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�  Z          \  [   X  O    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   W   Y   �     �	else if ((sprite_row + 195 < pixel_row) && (pixel_row < sprite_row + 201) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 81)) || ((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 180 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 230 < pixel_column) && (pixel_column < sprite_column + 241))))5�_�   i   k       l   j   I   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     0	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 1)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 220 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�   j               k   I   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   H   J   �     2	else if ((sprite_row + 160 < pixel_row) && (pixel_row < sprite_row + 171) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 70 < pixel_column) && (pixel_column < sprite_column + 131)) || ((sprite_column + 140 < pixel_column) && (pixel_column < sprite_column + 151)) || ((sprite_column + 200 < pixel_column) && (pixel_column < sprite_column + 211)) ||  ((sprite_column + 220 < pixel_column) && (pixel_column < sprite_column + 231)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�                    9        ����                                                                                                                                                                                                                                                                                                                                                             d     �   9   :   �    �   8   :   �      		// Row 51 - 90  �    else if ((sprite_row + 50 < pixel_row) && (pixel_row < sprite_row + 91) && (((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 210 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))           begin   !            winner_pix = 4'b1111;           end   	// Row 91 - 100  C    else if ((sprite_row + 90 < pixel_row) && (pixel_row < sprite_row + 101) && (((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 210 < pixel_column) && (pixel_column < sprite_column + 281))))           begin   !            winner_pix = 4'b1111;           end   // Row 51 - 1005�_�                     8        ����                                                                                                                                                                                                                                                                                                                                                             d�     �   8   9   �    �   7   9   �       	// Row 51 - 90  �    else if ((sprite_row + 50 < pixel_row) && (pixel_row < sprite_row + 91) && (((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 121)) || ((sprite_column + 170 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 210 < pixel_column) && (pixel_column < sprite_column + 221)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 281))))           begin   !            winner_pix = 4'b1111;           end   	// Row 91 - 100  C    else if ((sprite_row + 90 < pixel_row) && (pixel_row < sprite_row + 101) && (((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 51)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 181)) || ((sprite_column + 210 < pixel_column) && (pixel_column < sprite_column + 281))))           begin   !            winner_pix = 4'b1111;           end   
       end5��