Vim�UnDo� :$�t��?_AŞ@^���_(4"����1���   =   logic   [11:0]      alien2_row;            e       e   e   e    d	��    _�                             ����                                                                                                                                                                                                                                                                                                                                                             d	�D     �                   5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d	�J     �          /       5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d	�M     �          5       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d	�{     �          6      @// SV Module to Display One Copy of Alien A Through the VGA Port5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d	�}     �          6      @// SV Module to display One Copy of Alien A Through the VGA Port5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d	�     �          6      @// SV Module to display one Copy of Alien A Through the VGA Port5�_�                       %    ����                                                                                                                                                                                                                                                                                                                                                             d	��     �          6      @// SV Module to display one copy of Alien A Through the VGA Port5�_�      	                 *    ����                                                                                                                                                                                                                                                                                                                                                             d	��     �          6      @// SV Module to display one copy of alien A Through the VGA Port5�_�      
           	      )    ����                                                                                                                                                                                                                                                                                                                                                             d	��     �          6      ?// SV Module to display one copy of alienA Through the VGA Port5�_�   	              
      -    ����                                                                                                                                                                                                                                                                                                                                                             d	��     �          6      @// SV Module to display one copy of alien_A Through the VGA Port5�_�   
                    =    ����                                                                                                                                                                                                                                                                                                                                                             d	��     �          6      @// SV Module to display one copy of alien_A through the VGA Port5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d	��     �         6      // Module include 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d	��     �         8      @// addresses.  Future Updates will include automated motion for 5�_�                       0    ����                                                                                                                                                                                                                                                                                                                                                             d	�     �         8      E// addresses.  Future improvements will include automated motion for 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d	�     �         9      %// to implement automated motion for    	the Alien�         9      // the Alien5�_�                       .    ����                                                                                                                                                                                                                                                                                                                                                             d	�     �         8      .// to implement automated motion for the Alien5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d	�1     �         :      (// Created by Alexander Maso Winter 20235�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d	�;     �      C   :       5�_�                    	        ����                                                                                                                                                                                                                                                                                                                                                             d	�{     �      	           5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                             d	�}     �      
   s      *       input wire            vga_fast_clk,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d	�U     �      	   s      module alien_a(5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             d	��     �                	input  wire   [11:0]  btn_row,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d	��     �                	input  wire   [11:0]  btn_col5�_�                   %        ����                                                                                                                                                                                                                                                                                                                                                             d	��     �   $   %          logic [11:0]        btn_row_ff;5�_�                    %        ����                                                                                                                                                                                                                                                                                                                                                             d	��     �   $   %          logic [11:0]        btn_col_ff;5�_�                    $        ����                                                                                                                                                                                                                                                                                                                                                             d	��     �   #   $          // Internal ffs for Buttons5�_�                    )        ����                                                                                                                                                                                                                                                                                                                                                             d	��     �   (   )          btn_row_ff = 0;5�_�                    )        ����                                                                                                                                                                                                                                                                                                                                                             d	��     �   (   )          btn_col_ff = 0;5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �      
   l      '    input wire            vga_fast_clk,5�_�      !               	       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �      
   l      &    input wire            ga_fast_clk,5�_�       "           !   	       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �      
   l      %    input wire            a_fast_clk,5�_�   !   #           "   	       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �      
   l      $    input wire            _fast_clk,5�_�   "   $           #   	       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �      
   l      #    input wire            fast_clk,5�_�   #   %           $   	       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �      
   l      "    input wire            ast_clk,5�_�   $   &           %   	       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �      
   l      !    input wire            st_clk,5�_�   %   '           &   	       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �      
   l           input wire            t_clk,5�_�   &   (           '   	       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �      
   l          input wire            _clk,5�_�   '   )           (   
       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �   	      l      $    input wire            vga_rst_i,5�_�   (   *           )   
       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �   	      l      #    input wire            ga_rst_i,5�_�   )   +           *   
       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �   	      l      "    input wire            a_rst_i,5�_�   *   ,           +   
       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �   	      l      !    input wire            _rst_i,5�_�   +   -           ,          ����                                                                                                                                                                                                                                                                                                                                                             d	�     �   
                  output wire   [3:0]   vga_r,5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                                                             d	�     �   
             	output wire   [3:0]   vga_g,5�_�   -   /           .          ����                                                                                                                                                                                                                                                                                                                                                             d	�     �   
             	output wire   [3:0]   vga_b,5�_�   .   0           /          ����                                                                                                                                                                                                                                                                                                                                                             d	�     �   
             	output wire		      vga_hs,5�_�   /   1           0   
       ����                                                                                                                                                                                                                                                                                                                                                             d	�     �   
      h    �   
      h    5�_�   0   2           1          ����                                                                                                                                                                                                                                                                                                                                                             d	�      �   
      i           input wire            rst_i,5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                                                             d	�'     �         i      	output wire			  vga_vs,5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                                             d	�:     �         i      	output wire			  alien2_pix,5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                                                             d	�A     �   
      i          input wire            en,5�_�   4   6           5          ����                                                                                                                                                                                                                                                                                                                                                             d	�D     �         i      #	output wire  [3:0]			  alien2_pix,5�_�   5   7           6           ����                                                                                                                                                                                                                                                                                                                                                             d	�H     �   
      i      $    input wire                   en,5�_�   6   8           7   
       ����                                                                                                                                                                                                                                                                                                                                                             d	�K     �   	      i           input wire            rst_i,5�_�   7   9           8          ����                                                                                                                                                                                                                                                                                                                                                             d	�M     �   
      i           input wire               en,5�_�   8   :           9   	       ����                                                                                                                                                                                                                                                                                                                                                             d	�N     �      
   i          input wire            clk,5�_�   9   ;           :          ����                                                                                                                                                                                                                                                                                                                                                             d	�P     �   
      i          input wire              en,5�_�   :   <           ;           ����                                                                                                                                                                                                                                                                                                                                                             d	�[     �                reg  [3:0]      vga_r_reg;5�_�   ;   =           <           ����                                                                                                                                                                                                                                                                                                                                                             d	�[     �                reg  [3:0]      vga_g_reg;5�_�   <   >           =           ����                                                                                                                                                                                                                                                                                                                                                             d	�\     �                reg  [3:0]      vga_b_reg;5�_�   =   ?           >   
        ����                                                                                                                                                                                                                                                                                                                                                             d	�_     �   	      f      "    input wire              rst_i,5�_�   >   @           ?          ����                                                                                                                                                                                                                                                                                                                                                             d	�h     �         f      logic           vga_31_5_clk;5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                             d	�m     �                wire [31:0]     pix_num;   wire [3:0]      doutb;   logic           video_on;   logic [3:0]     vga_output;   lod4gic           vga_31_5_clk;5�_�   @   B           A           ����                                                                                                                                                                                                                                                                                                                                                             d	�n     �                &// Internals for VGA and ROM/RAM image5�_�   A   C           B           ����                                                                                                                                                                                                                                                                                                                                                             d	�y     �                // Internals for Ship   logic [11:0]        pixel_row;   !logic [11:0]        pixel_column;   logic [11:0]        ship_row;    logic [11:0]        ship_column;5�_�   B   D           C           ����                                                                                                                                                                                                                                                                                                                                                             d	��     �                video_on = 0;5�_�   C   E           D           ����                                                                                                                                                                                                                                                                                                                                                             d	��     �         Z      vga_output = 0;5�_�   D   F           E           ����                                                                                                                                                                                                                                                                                                                                                             d	��     �         Z      = 0;5�_�   E   G           F           ����                                                                                                                                                                                                                                                                                                                                                             d	��     �         Z       5�_�   F   I           G           ����                                                                                                                                                                                                                                                                                                                                                             d	��     �          [       5�_�   G   J   H       I   !        ����                                                                                                                                                                                                                                                                                                                                                             d	��     �       !       	   	.clock    	   (vga_31_5_clk),   	.rst	  	   (vga_rst_i),   	.video_on 	   (video_on),   	.horiz_sync	   (vga_hs),   	.vert_sync	   (vga_vs),   	.pixel_row     (pixel_row),   	.pixel_column  (pixel_column),   	.pix_num	   (pix_num)   );5�_�   I   K           J            ����                                                                                                                                                                                                                                                                                                                                                             d	��     �                 dtg dtg(5�_�   J   L           K            ����                                                                                                                                                                                                                                                                                                                                                             d	��     �                  5�_�   K   M           L            ����                                                                                                                                                                                                                                                                                                                                                             d	��     �                  5�_�   L   N           M            ����                                                                                                                                                                                                                                                                                                                                                             d	��     �                  5�_�   M   O           N   
        ����                                                                                                                                                                                                                                                                                                                                                             d	��     �   	      O      $//    input wire              rst_i,5�_�   N   P           O   
        ����                                                                                                                                                                                                                                                                                                                                                             d	��     �   	      O      #/    input wire              rst_i,5�_�   O   Q           P           ����                                                                                                                                                                                                                                                                                                                                                             d	��     �         O      enable = 0;5�_�   P   R           Q           ����                                                                                                                                                                                                                                                                                                                                                             d	��     �         O      = 0;5�_�   Q   S           R          ����                                                                                                                                                                                                                                                                                                                                                             d	�W     �         O      #	output wire  [3:0]	    alien2_pix,5�_�   R   T           S          ����                                                                                                                                                                                                                                                                                                                                                             d	�x     �         O      *	output wire  [63:0] [3:0]	    alien2_pix,5�_�   S   U           T           ����                                                                                                                                                                                                                                                                                                                                                             d	�     �         O       5�_�   T   V           U          ����                                                                                                                                                                                                                                                                                                                                                             d	��     �         P      // Internals5�_�   U   W           V          ����                                                                                                                                                                                                                                                                                                                                                             d	�     �         Q      :// Counter for pixel number: 6x6 Grid for Alien_2 = 64 pix5�_�   V   X           W           ����                                                                                                                                                                                                                                                                                                                                                             d	�     �         Q      :// Counter for pixel number: 8x6 Grid for Alien_2 = 64 pix5�_�   W   Y           X          ����                                                                                                                                                                                                                                                                                                                                                             d	�4     �         Q      alien2_pix = 0;5�_�   X   Z           Y   6       ����                                                                                                                                                                                                                                                                                                                                                             d	�P     �   5   6       
           end   -    // Row five through 10 of the ship sprite   �    else if (((ship_row + 4 < pixel_row) && (pixel_row < ship_row + 11)) && (ship_column < pixel_column) && (pixel_column < ship_column + 16))           begin   !            vga_output = 4'b1111;           end       else           begin   !            vga_output = 4'b0000;       end5�_�   Y   [           Z   ,       ����                                                                                                                                                                                                                                                                                                                                                             d	�S     �   +   ,       
           end       #    // Row three of the ship sprite   r    else if ((ship_row + 3 == pixel_row) && (ship_column + 2 < pixel_column) && (pixel_column < ship_column + 14))           begin   !            vga_output = 4'b1111;           end   "    // Row four of the ship sprite   r    else if ((ship_row + 4 == pixel_row) && (ship_column + 1 < pixel_column) && (pixel_column < ship_column + 15))           begin   !            vga_output = 4'b1111;5�_�   Z   \           [   &        ����                                                                                                                                                                                                                                                                                                                                                             d	�W     �   %   &          D    // ship is centered in the upper left corner | Row x Col / (0,0)5�_�   [   ]           \   '       ����                                                                                                                                                                                                                                                                                                                                                             d	�X     �   &   '          -    // Row one and Row two of the ship sprite5�_�   \   ^           ]   '       ����                                                                                                                                                                                                                                                                                                                                                             d	�Y     �   &   '          �    if (((ship_row < pixel_row) && (pixel_row < ship_row + 3)) && ((ship_column < (pixel_column + 6)) && (pixel_column < ship_column + 8)))5�_�   ]   _           ^   '       ����                                                                                                                                                                                                                                                                                                                                                             d	�Y     �   &   '                  begin5�_�   ^   `           _   '       ����                                                                                                                                                                                                                                                                                                                                                             d	�Z     �   &   '          !            vga_output = 4'b1111;5�_�   _   a           `   &        ����                                                                                                                                                                                                                                                                                                                                                             d	�\     �   %   *   9          5�_�   `   b           a          ����                                                                                                                                                                                                                                                                                                                                                             d	��     �         <           logic   [5:0]       counter;5�_�   a   c           b           ����                                                                                                                                                                                                                                                                                                                                                             d	��     �         <       5�_�   b   d           c          ����                                                                                                                                                                                                                                                                                                                                                             d	��     �         <    �         <    5�_�   c   e           d          ����                                                                                                                                                                                                                                                                                                                                                             d	��     �         =      logic   [11:0]      alien2_row;5�_�   d               e          ����                                                                                                                                                                                                                                                                                                                                                             d	��    �         =      logic   [11:0]      alien2_;5�_�   G           I   H   "        ����                                                                                                                                                                                                                                                                                                                                                             d	��     �   !   *        5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                             d	��     �      
   l          input wire            ,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             d	��     �              5��