Vim�UnDo� �k�J��r���;p|&��>FBP6�1A2  Y   !        if (sprite_column > 560)   ,                          dʛ    _�                     ,       ����                                                                                                                                                                                                                                                                                                                                                             dʚ    �  +  -  Y      !        if (sprite_column > 560) 5��