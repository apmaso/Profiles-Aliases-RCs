Vim�UnDo� 	�,lp6E޾��zg�r6<�Si���ːy;G   �                 �       �   �   �    d��    _�                             ����                                                                                                                                                                                                                                                                                                                                                             dhh     �                   5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             dh�     �         �      '	output wire    [3:0]	   alien2_output,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             dh�     �         �      module alien2(5�_�                       ,    ����                                                                                                                                                                                                                                                                                                                                                             dh�     �         �      '	output wire    [3:0]	   player_output,    �         �      ,    output wire                alien2_active5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             di     �         �      'logic   [11:0]              sprite_row;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             di     �         �      logic   [11:0]              ;5�_�                       #    ����                                                                                                                                                                                                                                                                                                                                                             di      �         �      *logic   [11:0]              sprite_column;5�_�      	                 "    ����                                                                                                                                                                                                                                                                                                                                                             di/     �         �      *logic   [11:0]              sprite_row_ff;5�_�      
           	      "    ����                                                                                                                                                                                                                                                                                                                                                             diO     �         �      -logic   [11:0]              sprite_column_ff;5�_�   	              
      "    ����                                                                                                                                                                                                                                                                                                                                                             diX     �         �      'logic   [3:0]               alien2_pix;5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                             diq     �         �    �         �    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             diu     �                'logic   [3:0]               player_pix;5�_�                       "    ����                                                                                                                                                                                                                                                                                                                                                             di~     �         �      ,logic   [11:0]              sprite_row_next;5�_�                          ����                                                                                                                                                                                                                                                                                                                                                           di�     �         �      &logic   [11:0]              _row_next;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                           di�     �         �      +logic   [11:0]             missle_row_next;5�_�                       "    ����                                                                                                                                                                                                                                                                                                                                                           di�     �         �      /logic   [11:0]              sprite_column_next;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                           di�     �                &logic                       move_left;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                           di�     �                )logic                       move_left_ff;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                           di�    �                +logic                       move_left_next;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                           dom     �                $logic                       active; 5�_�                            ����                                                                                                                                                                                                                                                                                                                                                           dos     �         �      *logic   [11:0]              missle_row_ff;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                           dou     �         �      -logic   [11:0]              missle_column_ff;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                           dov     �         �      ,logic   [11:0]              missle_row_next;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                           dow     �         �      /logic   [11:0]              missle_column_next;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                           dox     �         �      +logic   [23:0]              motion_counter;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                           do�     �          �          active = 1'b0;5�_�                        
    ����                                                                                                                                                                                                                                                                                                                                                           do�     �      !   �          alien2_pix = 4'b0000;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                           do�     �                    actidve = 1'b0;5�_�                    "       ����                                                                                                                                                                                                                                                                                                                                                           do�     �   !   "              sprite_column_ff = 312;5�_�                     "       ����                                                                                                                                                                                                                                                                                                                                                           do�     �   !   "              sprite_row_ff = 20;5�_�      !               "       ����                                                                                                                                                                                                                                                                                                                                                           do�     �   !   "              sprite_column = 312;5�_�       "           !   "       ����                                                                                                                                                                                                                                                                                                                                                           do�     �   !   "              sprite_row = 20;5�_�   !   #           "   "       ����                                                                                                                                                                                                                                                                                                                                                           do�     �   !   "              motion_counter = 0;5�_�   "   $           #   "       ����                                                                                                                                                                                                                                                                                                                                                           do�     �   !   "              move_left = 1'b0;5�_�   #   %           $   "        ����                                                                                                                                                                                                                                                                                                                                                           dp	     �   !   $   �      end5�_�   $   &           %   "        ����                                                                                                                                                                                                                                                                                                                                                           dp     �   !   #   �       5�_�   %   '           &   "       ����                                                                                                                                                                                                                                                                                                                                                           dp     �   "   $   �    �   "   #   �    5�_�   &   (           '   "       ����                                                                                                                                                                                                                                                                                                                                                           dp     �   "   $   �    �   "   #   �    5�_�   '   )           (   "       ����                                                                                                                                                                                                                                                                                                                                                           dp     �   !   "              5�_�   (   *           )   "       ����                                                                                                                                                                                                                                                                                                                                                           dp      �   !   #   �          player_pix = 4'b0000;5�_�   )   +           *   #       ����                                                                                                                                                                                                                                                                                                                                                           dp#     �   "   $   �          player_pix = 4'b0000;5�_�   *   ,           +           ����                                                                                                                                                                                                                                                                                                                                                           dp;     �      !   �      M    // Initializing Alien2 20 rows from the top of the screen. Rows 21 <-> 365�_�   +   -           ,       /    ����                                                                                                                                                                                                                                                                                                                                                           dp�     �      !   �      M    // Initializing Player 20 rows from the top of the screen. Rows 21 <-> 365�_�   ,   .           -       I    ����                                                                                                                                                                                                                                                                                                                                                           dp�     �      !   �      P    // Initializing Player 20 rows from the bottom of the screen. Rows 21 <-> 365�_�   -   /           .       Q    ����                                                                                                                                                                                                                                                                                                                                                           dp�     �      !   �      Q    // Initializing Player 20 rows from the bottom of the screen. Rows 451 <-> 365�_�   .   0           /   "       ����                                                                                                                                                                                                                                                                                                                                                           dp�     �   !   #   �          player_row = 4'b0000;5�_�   /   1           0   !   6    ����                                                                                                                                                                                                                                                                                                                                                           dp�     �       "   �      >    // and close to centered as possible. Columns: 313 <-> 3285�_�   0   2           1   !   >    ����                                                                                                                                                                                                                                                                                                                                                           dp�     �       "   �      >    // and close to centered as possible. Columns: 311 <-> 3285�_�   1   3           2   !   =    ����                                                                                                                                                                                                                                                                                                                                                           dp�     �       "   �      >    // and close to centered as possible. Columns: 311 <-> 3355�_�   2   4           3   !   6    ����                                                                                                                                                                                                                                                                                                                                                           dp�     �       "   �      >    // and close to centered as possible. Columns: 311 <-> 3255�_�   3   5           4   !   >    ����                                                                                                                                                                                                                                                                                                                                                           dp�     �       "   �      >    // and close to centered as possible. Columns: 313 <-> 3255�_�   4   6           5   !   6    ����                                                                                                                                                                                                                                                                                                                                                           dq     �       "   �      >    // and close to centered as possible. Columns: 313 <-> 3255�_�   5   7           6   !   6    ����                                                                                                                                                                                                                                                                                                                                                           drW     �       "   �      >    // and close to centered as possible. Columns: 311 <-> 3255�_�   6   8           7   !   >    ����                                                                                                                                                                                                                                                                                                                                                           dr\     �       "   �      >    // and close to centered as possible. Columns: 313 <-> 3255�_�   7   9           8   #       ����                                                                                                                                                                                                                                                                                                                                                           dr`     �   "   $   �          player_column = 4'b0000;5�_�   8   :           9   ,       ����                                                                                                                                                                                                                                                                                                                                                           drn     �   +   -   �      �    active = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 17));5�_�   9   ;           :   ,   =    ����                                                                                                                                                                                                                                                                                                                                                           drx     �   +   -   �      �    active = ((player_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 17));5�_�   :   <           ;   ,   F    ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   +   -   �      �    active = ((player_row < pixel_row) && (pixel_row < player_row + 17) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 17));5�_�   ;   =           <   ,   Q    ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   +   -   �      �    active = ((player_row < pixel_row) && (pixel_row < player_row + 11) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 17));5�_�   <   >           =   ,   M    ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   +   -   �      �    active = ((player_row < pixel_row) && (pixel_row < player_row + 11) && (e_column < pixel_column) && (pixel_column < sprite_column + 17));5�_�   =   ?           >   ,   �    ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   +   -   �      �    active = ((player_row < pixel_row) && (pixel_row < player_row + 11) && (player_column < pixel_column) && (pixel_column < sprite_column + 17));5�_�   >   @           ?   ,   �    ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   +   -   �      �    active = ((player_row < pixel_row) && (pixel_row < player_row + 11) && (player_column < pixel_column) && (pixel_column < player_column + 17));5�_�   ?   A           @   /       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   .   0   �      P    // Sprite data for Alien2....  I can make this logic much simpler, if needed5�_�   @   B           A   0        ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          +    // Row one & two of Alien2's Sprite    5�_�   A   C           B   0        ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row  + 3) && (sprite_column + 6 < pixel_column) && (pixel_column < sprite_column + 11))5�_�   B   D           C   0        ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  begin5�_�   C   E           D   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          !            alien2_pix = 4'b1111;5�_�   D   F           E   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  end   5�_�   E   G           F   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          #    // Row 3 & 4 of Alien2's Sprite5�_�   F   H           G   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          �    else if ((sprite_row + 2 < pixel_row) && (pixel_row < sprite_row  + 5) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 13))5�_�   G   I           H   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  begin5�_�   H   J           I   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          !            alien2_pix = 4'b1111;5�_�   I   K           J   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  end   5�_�   J   L           K   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          #    // Row 5 & 6 of Alien2's Sprite5�_�   K   M           L   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          �    else if ((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 7) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 15))5�_�   L   N           M   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  begin5�_�   M   O           N   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          !            alien2_pix = 4'b1111;5�_�   N   P           O   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  end5�_�   O   Q           P   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          #    // Row 7 & 8 of Alien2's Sprite5�_�   P   R           Q   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          �    else if ((sprite_row + 6 < pixel_row) && (pixel_row < sprite_row  +  9) && (pixel_column != sprite_column + 5) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 11) && (pixel_column != sprite_column + 12))5�_�   Q   S           R   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  begin5�_�   R   T           S   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          !            alien2_pix = 4'b1111;5�_�   S   U           T   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  end5�_�   T   V           U   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          $    // Row 9 & 10 of Alien2's Sprite5�_�   U   W           V   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          �    else if ((sprite_row + 8 < pixel_row) && (pixel_row < sprite_row + 11) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 17))5�_�   V   X           W   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  begin5�_�   W   Y           X   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          !            alien2_pix = 4'b1111;5�_�   X   Z           Y   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  end5�_�   Y   [           Z   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          %    // Row 11 & 12 of Alien2's Sprite5�_�   Z   \           [   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          �    else if ((sprite_row + 10 < pixel_row) && (pixel_row < sprite_row  + 13) && ((sprite_column + 5 == pixel_column) || (sprite_column + 6 == pixel_column) || (pixel_column == sprite_column + 11) || (pixel_column == sprite_column + 12)))5�_�   [   ]           \   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  begin5�_�   \   ^           ]   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          !            alien2_pix = 4'b1111;5�_�   ]   _           ^   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  end5�_�   ^   `           _   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          %    // Row 13 & 14 of Alien2's Sprite5�_�   _   a           `   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0         �    else if ((sprite_row + 12 < pixel_row) && (pixel_row < sprite_row  + 15) && (pixel_column != sprite_column + 1) && (pixel_column != sprite_column + 2) && (pixel_column != sprite_column + 5) && (pixel_column != sprite_column + 6) && (pixel_column != sprite_column + 11) && (pixel_column != sprite_column + 12) && (pixel_column != sprite_column + 15) && (pixel_column != sprite_column + 16))5�_�   `   b           a   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  begin5�_�   a   c           b   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          !            alien2_pix = 4'b1111;5�_�   b   d           c   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  end5�_�   c   e           d   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          %    // Row 15 & 16 of Alien2's Sprite5�_�   d   f           e   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0         �    else if ((sprite_row + 14 < pixel_row) && (pixel_row < sprite_row  + 17) && (pixel_column == sprite_column + 1) && (pixel_column == sprite_column + 2) && (pixel_column == sprite_column + 5) && (pixel_column == sprite_column + 6) && (pixel_column == sprite_column + 11) && (pixel_column == sprite_column + 12) && (pixel_column == sprite_column + 15) && (pixel_column == sprite_column + 16))5�_�   e   g           f   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  begin5�_�   f   h           g   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          !            alien2_pix = 4'b1111;5�_�   g   i           h   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  end 5�_�   h   j           i   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0              else5�_�   i   k           j   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  begin5�_�   j   l           k   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          !            alien2_pix = 4'b0000;5�_�   k   m           l   0       ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0                  end5�_�   l   n           m   0        ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   0          end5�_�   m   o           n   0        ����                                                                                                                                                                                                                                                                                                                                                           dr�     �   /   3   q       5�_�   n   p           o   0        ����                                                                                                                                                                                                                                                                                                                                                           ds3     �   /   H   s       5�_�   o   q           p   0       ����                                                                                                                                                                                                                                                                                                                                                           ds@     �   /   1   �      =        // Row one and two of the player's sprite            5�_�   p   r           q   1        ����                                                                                                                                                                                                                                                                                                                                                           dsr     �   ?   A          �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 11)) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 16))�   :   <          x    else if ((sprite_row + 4 == pixel_row) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 15))�   5   7          x    else if ((sprite_row + 3 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 14))�   0   2          i    if ((sprite_row < pixel_row) && (pixel_row < sprite_row  + 3) && (pixel_column == sprite_column + 8))5�_�   q   s           r   1        ����                                                                                                                                                                                                                                                                                                                                                           ds�     �   ?   A          �    else if (((player_row + 4 < pixel_row) && (pixel_row < player_row  + 11)) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 16))�   :   <          x    else if ((player_row + 4 == pixel_row) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 15))�   5   7          x    else if ((player_row + 3 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 14))�   0   2          i    if ((player_row < pixel_row) && (pixel_row < player_row  + 3) && (pixel_column == sprite_column + 8))5�_�   r   t           s   3        ����                                                                                                                                                                                                                                                                                                                                                           ds�     �   E   G                      vga_output = doutb;�   A   C          !            vga_output = 4'b1111;�   <   >          !            vga_output = 4'b1111;�   7   9          !            vga_output = 4'b1111;�   2   4          !            vga_output = 4'b1111;5�_�   s   u           t   F       ����                                                                                                                                                                                                                                                                                                                                                           ds�     �   E   G   �                  player_pix = doutb;5�_�   t   v           u   F       ����                                                                                                                                                                                                                                                                                                                                                           ds�     �   E   G   �                  player_pix = ;5�_�   u   w           v   I       ����                                                                                                                                                                                                                                                                                                                                                           dt     �   H   K   �             5�_�   v   x           w   H        ����                                                                                                                                                                                                                                                                                                                                                           dt     �   F   H   �              end    �   G   I   �       5�_�   w   y           x   �       ����                                                                                                                                                                                                                                                                                                                                                           dtu     �   �   �   �      "assign alien2_output = alien2_pix;5�_�   x   z           y   �       ����                                                                                                                                                                                                                                                                                                                                                           dtz     �   �   �   �      assign alien2_active = active; 5�_�   y   {           z   �       ����                                                                                                                                                                                                                                                                                                                                                           dt�     �   �   �   �      assign player_active = active; 5�_�   z   |           {   �       ����                                                                                                                                                                                                                                                                                                                                                           dt�     �   �   �   �      assign player_enable = active; 5�_�   {   }           |   �       ����                                                                                                                                                                                                                                                                                                                                                           dt�     �   �   �   �      "assign player_output = alien2_pix;5�_�   |   ~           }   �        ����                                                                                                                                                                                                                                                                                                                                                           dt�     �   �   �           assign move_left = move_left_ff;5�_�   }   �           ~   �        ����                                                                                                                                                                                                                                                                                                                                                           dt�     �   �   �          "assign sprite_row = sprite_row_ff;5�_�   ~   �          �   �        ����                                                                                                                                                                                                                                                                                                                                                           dt�     �   �   �          (assign sprite_column = sprite_column_ff;5�_�   �   �   �       �          ����                                                                                                                                                                                                                                                                                                                                                           dt�     �         �    �         �    5�_�   �   �           �      $    ����                                                                                                                                                                                                                                                                                                                                                           dt�     �         �      8    input  wire    [11:0]      pixel_row, pixel_column, 5�_�   �   �           �      -    ����                                                                                                                                                                                                                                                                                                                                                           dt�     �         �      6    input  wire    [11:0]      btn_row, pixel_column, 5�_�   �   �           �      2    ����                                                                                                                                                                                                                                                                                                                                                           dt�     �         �      4    input  wire    [11:0]      btn_row, btn_column, 5�_�   �   �           �   K   S    ����                                                                                                                                                                                                                                                                                                                                                           duf     �   J   M   �      S// Additional combinational block for FSM used in implemention of motion for Alien25�_�   �   �           �   r        ����                                                                                                                                                                                                                                                                                                                                                           duw     �   q   t   �       5�_�   �   �           �   r        ����                                                                                                                                                                                                                                                                                                                                                           duy     �   q   s   �       5�_�   �   �           �   r       ����                                                                                                                                                                                                                                                                                                                                                           du�     �   q   s   �      */5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                                                           du�     �   �   �   �       5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                                                           du�     �   J   L   �      S// Additional combinational block for FSM used in implemention of motion of Missles5�_�   �   �           �   K   R    ����                                                                                                                                                                                                                                                                                                                                                           du�     �   J   M   �      R// Additional comb and ff  block for FSM used in implemention of motion of Missles5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                                                           du�     �   J   L   �      G// Additional comb and ff  block for FSM used in implemention of motion5�_�   �   �           �   L   &    ����                                                                                                                                                                                                                                                                                                                                                           du�     �   K   N   �      &// Do not need this yet, first moving 5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                                                           dv     �   �   �   �       5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                           dv"     �   �   �   �    �   �   �   �    5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                           dv&     �   �   �   �      assign player_column = btn_col;5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                           dv+     �   �   �   �      assign player_column = btn_row;5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                           dv-     �   �   �   �      assign player_= btn_row;5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                           dv8     �   �   �   �      assign player_enable = enalbe; 5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                           dv;     �   �   �   �       assign player_enable = enaxlbe; 5�_�   �   �           �   �       ����                                                                                                                                                                                                                                                                                                                                                           dv=     �   �   �   �      assign player_enable = enabe; 5�_�   �   �           �   -   
    ����                                                                                                                                                                                                                                                                                                                                                           dvG     �   ,   .   �      �    active = ((player_row < pixel_row) && (pixel_row < player_row + 11) && (player_column < pixel_column) && (pixel_column < player_column + 16));5�_�   �   �           �   �        ����                                                                                                                                                                                                                                                                                                                                                           dv�     �   �   �          assign player_enable = enable; 5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                                                           dw     �   ,   .   �      �    enable = ((player_row < pixel_row) && (pixel_row < player_row + 11) && (player_column < pixel_column) && (pixel_column < player_column + 16));5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                           dw     �         �      &	output wire    [3:0]	   player_output5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                           dw     �         �      	i5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                           dw"     �         �    �         �    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                           dw$     �                	5�_�   �   �           �      /    ����                                                                                                                                                                                                                                                                                                                                                           dw'     �         �      1    input  wire    [11:0]      btn_row, btn_col, 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                           dw/     �         �      .    input  wire    [11:0]      player_enable, 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                           dw8     �         �      .    output wire    [11:0]      player_enable, 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                           dw>     �         �      .    output wire    [11:0]      player_enable, 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                           dwB    �         �      )    output wire           player_enable, 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                           d��     �         �      1    input  wire    [11:0]      btn_row, btn_col, 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                           d��     �         �      *    input  wire    [11:0]      , btn_col, 5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                           d��     �         �      )    input  wire    [11:0]       btn_col, 5�_�   �               �   �        ����                                                                                                                                                                                                                                                                                                                                                           d��    �   �   �          assign player_row = btn_row;5�_�   �       �   �   �          ����                                                                                                                                                                                                                                                                                                                                                           dt�     �         �    �         �      8    input  wire    [11:0]      pixel_row, pixel_column,    &	output wire    [3:0]	   player_output5�_�   �           �   �          ����                                                                                                                                                                                                                                                                                                                                                           dt�     �         �    �         �      8    input  wire    [11:0]      pixel_row, pixel_column,    &	output wire    [3:0]	   player_output5�_�   ~           �      �        ����                                                                                                                                                                                                                                                                                                                                                           dt�     �   �   �        5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             di�     �         �    �         �      6logic   [11:0]              _missle_column_ffrow_next;5��