Vim�UnDo� L�p }�q#)����-�FR��m"�5 ��   �       sprite_column = 400;   #                      d�    _�                     -       ����                                                                                                                                                                                                                                                                                                                                                             d�}     �   ,   .   �      �     active2 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 61));    5�_�                    /       ����                                                                                                                                                                                                                                                                                                                                                             d�     �   .   0   �      �     active3 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 101));5�_�                    1       ����                                                                                                                                                                                                                                                                                                                                                             d��     �   0   2   �      �     active4 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 141));5�_�                    +   �    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   *   ,   �      �    active1 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 21));5�_�                    -   ]    ����                                                                                                                                                                                                                                                                                                                                                             d�)     �   ,   .   �      �    active2 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 61));    5�_�                    -   �    ����                                                                                                                                                                                                                                                                                                                                                             d�.     �   ,   .   �      �    active2 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 61));    5�_�                    /   _    ����                                                                                                                                                                                                                                                                                                                                                             d�5     �   .   0   �      �    active3 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 101));5�_�      	              /   �    ����                                                                                                                                                                                                                                                                                                                                                             d�:     �   .   0   �      �    active3 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 101));5�_�      
           	   1   �    ����                                                                                                                                                                                                                                                                                                                                                             d�@     �   0   2   �      �    active4 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 141));5�_�   	              
   1   _    ����                                                                                                                                                                                                                                                                                                                                                             d�G     �   0   2   �      �    active4 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 281));5�_�   
                 +   G    ����                                                                                                                                                                                                                                                                                                                                                             d�U     �   *   ,   �      �    active1 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 41));5�_�                    -   G    ����                                                                                                                                                                                                                                                                                                                                                             d�W     �   ,   .   �      �    active2 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 121));    5�_�                    /   G    ����                                                                                                                                                                                                                                                                                                                                                             d�X     �   .   0   �      �    active3 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 201));5�_�                    1   G    ����                                                                                                                                                                                                                                                                                                                                                             d�Z     �   0   2   �      �    active4 = ((sprite_row < pixel_row) && (pixel_row < sprite_row + 17) && (sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 281));5�_�                    (       ����                                                                                                                                                                                                                                                                                                                                                             d�d     �   '   )   �      <    // Barrier Sprite's are 16 rows by 20 columns of pixels 5�_�                    (   (    ����                                                                                                                                                                                                                                                                                                                                                             d�f     �   '   )   �      <    // Barrier Sprite's are 32 rows by 20 columns of pixels 5�_�                    )       ����                                                                                                                                                                                                                                                                                                                                                             d�l     �   (   *   �      W    // There are 20 pixels between each barrier sprite --> Offsets are multiples of 40 5�_�                    ,   $    ����                                                                                                                                                                                                                                                                                                                                                             d�u     �   +   -   �      &    // Second sprite --> Offset of 40 5�_�                    .   #    ����                                                                                                                                                                                                                                                                                                                                                             d�x     �   -   /   �      %    // Third sprite --> Offset of 80 5�_�                    0   $    ����                                                                                                                                                                                                                                                                                                                                                             d�z     �   /   1   �      %    // Fourth sprite --> Offset of 805�_�                    .   $    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   -   /   �      &    // Third sprite --> Offset of 120 5�_�                    0   #    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   /   1   �      $    // Fourth sprite --> Offset of 05�_�                    5   ;    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   4   6   �      t    if ((pixel_row == sprite_row  + 1) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 19))5�_�                    5   q    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   4   6   �      t    if ((pixel_row == sprite_row  + 1) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 19))5�_�                    5   p    ����                                                                                                                                                                                                                                                                                                                                                             d��    �   4   6   �      t    if ((pixel_row == sprite_row  + 1) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 17))5�_�                    :   ?    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   9   ;   �      x    else if ((sprite_row + 2 == pixel_row) && (sprite_column + 1 < pixel_column) && (pixel_column < sprite_column + 20))5�_�                    :   t    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   9   ;   �      x    else if ((sprite_row + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 20))5�_�                    :   u    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   9   ;   �      x    else if ((sprite_row + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 30))5�_�                    ?   �    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   >   @   �      �    else if ((sprite_row + 2 < pixel_row) && (pixel_row < sprite_row  + 10) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 21))5�_�                    5       ����                                                                                                                                                                                                                                                                                                                            5   &       5          v       d��     �   4   6   �      t    if ((pixel_row == sprite_row  + 1) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�                     5       ����                                                                                                                                                                                                                                                                                                                            5   &       5          v       d��     �   4   6   �      s    if ((pixel_row = sprite_row  + 1) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�      !               5       ����                                                                                                                                                                                                                                                                                                                            5   &       5          v       d��     �   4   6   �      r    if ((pixel_row  sprite_row  + 1) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�       "           !   5   #    ����                                                                                                                                                                                                                                                                                                                            5   &       5          v       d��     �   4   6   �      s    if ((pixel_row < sprite_row  + 1) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   !   #           "   5   &    ����                                                                                                                                                                                                                                                                                                                            5   &       5          v       d��     �   4   6   �      u    if ((pixel_row < sprite_row  + xx1) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   "   $           #   5   	    ����                                                                                                                                                                                                                                                                                                                            5   &       5          v       d��     �   4   6   �      a    if ((pixel_row) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   #   %           $   5   	    ����                                                                                                                                                                                                                                                                                                                            5   &       5          v       d��     �   4   6   �      c    if ((< pixel_row) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   $   &           %   5   $    ����                                                                                                                                                                                                                                                                                                                            5   &       5          v       d�     �   4   6   �      n    if ((sprite_row < pixel_row) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   %   '           &   5   $    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      n    if ((sprite_row < pixel_row) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))�   5   6   �    5�_�   &   (           '   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      �    if ((sprite_row < pixel_row) && ((sprite_row < pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   '   )           (   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      �    if ((sprite_row < pixel_row) && (sprite_row < pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   (   *           )   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      �    if ((sprite_row < pixel_row) && (prite_row < pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   )   +           *   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      �    if ((sprite_row < pixel_row) && (rite_row < pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   *   ,           +   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      �    if ((sprite_row < pixel_row) && (ite_row < pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   +   -           ,   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      �    if ((sprite_row < pixel_row) && (te_row < pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   ,   .           -   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      �    if ((sprite_row < pixel_row) && (e_row < pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   -   /           .   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      �    if ((sprite_row < pixel_row) && (_row < pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   .   0           /   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �          if ((sprite_row < pixel_row) && (row < pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   /   1           0   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      ~    if ((sprite_row < pixel_row) && (ow < pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   0   2           1   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      }    if ((sprite_row < pixel_row) && (w < pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   1   3           2   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      |    if ((sprite_row < pixel_row) && ( < pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   2   4           3   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      {    if ((sprite_row < pixel_row) && (< pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   3   5           4   5   %    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      z    if ((sprite_row < pixel_row) && ( pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   4   6           5   5   .    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�     �   4   6   �      y    if ((sprite_row < pixel_row) && (pixel_row) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   5   7           6   4       ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�%     �   3   5   �      '    // Row one of Barrier1's Sprite    5�_�   6   8           7   4       ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�+     �   3   5   �      '    // Row 1&2 of Barrier1's Sprite    5�_�   7   9           8   4       ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�+     �   3   5   �      (    // Row 1 &2 of Barrier1's Sprite    5�_�   8   :           9   5   A    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�6     �   4   6   �      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   9   ;           :   5   C    ����                                                                                                                                                                                                                                                                                                                            5           5          v       d�8     �   4   6   �      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) &&(sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   :   <           ;   :       ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�Q     �   9   ;   �      x    else if ((sprite_row + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))�   :   ;   �    5�_�   ;   =           <   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�T     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) sprite_row + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   <   >           =   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�T     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)sprite_row + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   =   ?           >   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�T     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)prite_row + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   >   @           ?   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�U     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)rite_row + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   ?   A           @   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�U     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)ite_row + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   @   B           A   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�U     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)te_row + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   A   C           B   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�U     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)e_row + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   B   D           C   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�U     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)_row + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   C   E           D   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�U     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)row + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   D   F           E   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�U     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)ow + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   E   G           F   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�U     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)w + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   F   H           G   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�U     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) + 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   G   I           H   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�U     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)+ 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   H   J           I   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�U     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) 2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   I   K           J   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�U     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)2 == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   J   L           K   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�V     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) == pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   K   M           L   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�V     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)== pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   L   N           M   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�V     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)= pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   M   O           N   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�V     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   N   P           O   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�V     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)pixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   O   Q           P   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�V     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)ixel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   P   R           Q   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�W     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)xel_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   Q   S           R   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�W     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)el_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   R   T           S   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�W     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)l_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   S   U           T   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�W     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)_row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   T   V           U   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�W     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)row) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   U   W           V   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�W     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)ow) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   V   X           W   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�X     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)w) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   W   Y           X   :   F    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�Y     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3)) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   X   Z           Y   :   D    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�[     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   Y   [           Z   :       ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�a     �   9   ;   �      �    else if (((sprite_row < pixel_row) && (pixel_row < sprite_row + 5) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   Z   \           [   :       ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�h     �   9   ;   �      �    else if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 5) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   [   ]           \   9       ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d�u     �   8   :   �          // Row 2 5�_�   \   ^           ]   >       ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d��     �   =   ?   �          // Rows 3 - 9 5�_�   ]   _           ^   >       ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d��     �   =   ?   �          // Rows 5 - 9 5�_�   ^   `           _   ?       ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d��     �   >   @   �      �    else if ((sprite_row + 2 < pixel_row) && (pixel_row < sprite_row  + 10) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 41))5�_�   _   a           `   ?   J    ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d��     �   >   @   �      �    else if ((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 10) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 41))5�_�   `   c           a   C       ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d��     �   B   D   �          // Row 105�_�   a   d   b       c   D       ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if ((sprite_row + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))�   D   E   �    5�_�   c   e           d   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �         else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) sprite_row + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   d   f           e   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �         else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)sprite_row + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   e   g           f   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �         else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)prite_row + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   f   h           g   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �         else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)rite_row + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   g   i           h   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �         else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)ite_row + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   h   j           i   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �         else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)te_row + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   i   k           j   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �         else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)e_row + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   j   l           k   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �          else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)_row + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   k   m           l   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)row + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   l   n           m   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)ow + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   m   o           n   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)w + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   n   p           o   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   o   q           p   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)+ 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   p   r           q   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   q   s           r   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   r   t           s   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)0 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   s   u           t   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   t   v           u   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)== pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   u   w           v   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)= pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   v   x           w   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   w   y           x   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   x   z           y   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)ixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   y   {           z   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)xel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   z   |           {   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)el_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   {   }           |   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)l_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   |   ~           }   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   }              ~   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   ~   �              D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)ow) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�      �           �   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)w) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   D   L    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19)) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   D       ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if (((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   D       ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if ((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   D   I    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row  + 19) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   D   I    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row  + 9) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   D   I    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row  + ) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   D   E    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d��     �   C   E   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row  + 21) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   D   �    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d�     �   C   E   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   D   �    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d�     �   C   E   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + )) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   D   �    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d�5     �   C   E   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 15)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   D   �    ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d�<     �   C   E   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 15)) || ((sprite_column + 26 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   H       ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d�D     �   G   I   �          // Row 11 5�_�   �   �           �   H       ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d�G     �   G   I   �          // Row 21 5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d�V     �   H   J   �      �    else if ((sprite_row + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))�   I   J   �    5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            ?          ?   K       v   K    d�Y     �   H   J   �      �    else if ((8sprite_row + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�c     �   H   J   �      �    else if ((sprite_row + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))�   I   J   �    5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�g     �   H   J   �         else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) sprite_row + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �         else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)sprite_row + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �         else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)prite_row + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �         else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)rite_row + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �         else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)ite_row + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �         else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)te_row + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �         else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)e_row + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �          else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)_row + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)row + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)ow + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)w + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) + 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)+ 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) 11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)11 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)1 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)== pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)= pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�h     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�i     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)ixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�i     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)xel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�i     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)el_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�i     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)l_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�i     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�i     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�i     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)ow) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�j     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)w) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   L    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�j     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21)) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�p     �   H   J   �      �    else if (((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�t     �   H   J   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�v     �   H   J   �      �    else if ((sprite_row + 28 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   I    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�{     �   H   J   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   �    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d��     �   H   J   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 7)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   �    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d��     �   H   J   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + )) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   �    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d��     �   H   J   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 13)) || ((sprite_column + 14 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   I   �    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d��     �   H   J   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 13)) || ((sprite_column + 28 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d��     �   L   N   �          // Rows 12 & 135�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d��     �   L   N   �          // Rows 23 & 135�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d��     �   L   N   �          // Rows 23 - 135�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d��     �   M   O   �      �    else if ((sprite_row + 11 < pixel_row) && (pixel_row < sprite_row + 14) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 6)) || ((sprite_column + 15 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   N   J    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d��     �   M   O   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 14) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 6)) || ((sprite_column + 15 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   N   �    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�     �   M   O   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 6)) || ((sprite_column + 15 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   N   �    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�&     �   M   O   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 15 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   N   �    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�,     �   M   O   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 30 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   S   �    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�4     �   R   T   �      �    else if ((sprite_row + 13 < pixel_row) && (pixel_row < sprite_row + 17) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 5)) || ((sprite_column + 16 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�   �   �           �   S   �    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�E     �   R   T   �      �    else if ((sprite_row + 13 < pixel_row) && (pixel_row < sprite_row + 17) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 5)) || ((sprite_column + 16 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�   �   �           �   S   �    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�[     �   R   T   �      �    else if ((sprite_row + 13 < pixel_row) && (pixel_row < sprite_row + 17) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 5)) || ((sprite_column + 32 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�a     �   Q   S   �          // Row 14, 15 and 16 5�_�   �   �           �   S       ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�l     �   R   T   �      �    else if ((sprite_row + 13 < pixel_row) && (pixel_row < sprite_row + 17) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 9)) || ((sprite_column + 32 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�   �   �           �   S   J    ����                                                                                                                                                                                                                                                                                                                            D          D   K       v   K    d�p     �   R   T   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 17) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 9)) || ((sprite_column + 32 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�   �   �           �   Z        ����                                                                                                                                                                                                                                                                                                                            W           4           v        d£     �   Y   Z          z    else if ((pixel_row == sprite_row  + 1) && (sprite_column + 42 < pixel_column) && (pixel_column < sprite_column + 59))5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d£     �   Y   Z                  begin5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d£     �   Y   Z          "            barrier_pix = 4'b1111;5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¤     �   Y   Z                  end   5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¤     �   Y   Z              // Row 2 5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¤     �   Y   Z          y    else if ((sprite_row + 2 == pixel_row) && (sprite_column + 41 < pixel_column) && (pixel_column < sprite_column + 60))5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¤     �   Y   Z                  begin5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¥     �   Y   Z          "            barrier_pix = 4'b1111;5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¥     �   Y   Z                  end   5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¥     �   Y   Z              // Rows 3 - 9 5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¦     �   Y   Z          �    else if ((sprite_row + 2 < pixel_row) && (pixel_row < sprite_row  + 10) && (sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 61))5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¦     �   Y   Z                  begin5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¦     �   Y   Z          "            barrier_pix = 4'b1111;5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d§     �   Y   Z                  end5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d§     �   Y   Z              // Row 105�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d§     �   Y   Z          �    else if ((sprite_row + 10 == pixel_row) && (((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 48)) || ((sprite_column + 53 < pixel_column) && (pixel_column < sprite_column + 61))))5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d§     �   Y   Z                  begin5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¨     �   Y   Z          "            barrier_pix = 4'b1111;5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¨     �   Y   Z                  end5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d©     �   Y   Z              // Row 11 5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d©     �   Y   Z          �    else if ((sprite_row + 11 == pixel_row) && (((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 47)) || ((sprite_column + 54 < pixel_column) && (pixel_column < sprite_column + 61))))5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d©     �   Y   Z                  begin5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d©     �   Y   Z          "            barrier_pix = 4'b1111;5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        dª     �   Y   Z                  end5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        dª     �   Y   Z              // Rows 12 & 135�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        dª     �   Y   Z          �    else if ((sprite_row + 11 < pixel_row) && (pixel_row < sprite_row + 14) && (((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 46)) || ((sprite_column + 55 < pixel_column) && (pixel_column < sprite_column + 61))))5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d«     �   Y   Z                  begin5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d«     �   Y   Z          "            barrier_pix = 4'b1111;5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d«     �   Y   Z                  end5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¬     �   Y   Z              // Row 14, 15 and 16 5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¬     �   Y   Z          �    else if ((sprite_row + 13 < pixel_row) && (pixel_row < sprite_row + 17) && (((sprite_column + 40 < pixel_column) && (pixel_column < sprite_column + 45)) || ((sprite_column + 56 < pixel_column) && (pixel_column < sprite_column + 61))))5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d­     �   Y   Z                  begin5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d­     �   Y   Z          "            barrier_pix = 4'b1111;5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           4           v        d®     �   Y   Z                  end5�_�   �   �           �   Y   .    ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¶     �   X   Z   �      8    // Row one of Barrier2's Sprite (Offset = 40 pix)   5�_�   �   �           �   \   .    ����                                                                                                                                                                                                                                                                                                                            W           4           v        dº     �   [   ]   �      8    // Row one of Barrier3's Sprite (Offset = 80 pix)   5�_�   �   �           �   \   .    ����                                                                                                                                                                                                                                                                                                                            W           4           v        d»     �   [   ]   �      8    // Row one of Barrier3's Sprite (Offset = 10 pix)   5�_�   �   �           �   \   /    ����                                                                                                                                                                                                                                                                                                                            W           4           v        d¼     �   [   ]   �      8    // Row one of Barrier3's Sprite (Offset = 10 pix)   5�_�   �   �   �       �   Z        ����                                                                                                                                                                                                                                                                                                                            W           5           v        d��     �   Y   ~   �       �   Z   [   �    5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           5           v        d��     �   Y   [   �      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   �   �           �   Z       ����                                                                                                                                                                                                                                                                                                                            W           5           v        d��     �   Y   [   �      �    if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   �   �           �   X        ����                                                                                                                                                                                                                                                                                                                            W           5           v        d��     �   W   X           5�_�   �   �           �   X       ����                                                                                                                                                                                                                                                                                                                            W           5           v        d��     �   W   Y   �      8    // Row one of Barrier2's Sprite (Offset = 80 pix)   5�_�   �   �           �   Y   Z    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d��     �   X   Z   �      �    else if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) && (sprite_column + 4 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   �   �   �       �   Y   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�     �   X   Z   �      �    else if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) && (sprite_column + 84 < pixel_column) && (pixel_column < sprite_column + 37))5�_�   �   �           �   ^   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�*     �   ]   _   �      �    else if ((sprite_row + 2 < pixel_row) && (pixel_row < sprite_row + 5) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 39))5�_�   �   �           �   ^   ^    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�/     �   ]   _   �      �    else if ((sprite_row + 2 < pixel_row) && (pixel_row < sprite_row + 5) && (sprite_column + 2 < pixel_column) && (pixel_column < sprite_column + 119))5�_�   �   �           �   c   ^    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�7     �   b   d   �      �    else if ((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) && (sprite_column < pixel_column) && (pixel_column < sprite_column + 41))5�_�   �   �   �       �   c   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�S     �   b   d   �      �    else if ((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) && (sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 41))5�_�   �   �           �   h   `    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�[     �   g   i   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 15)) || ((sprite_column + 26 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�   �   �           �   h   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�a     �   g   i   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 15)) || ((sprite_column + 26 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�   �   �           �   h   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�d     �   g   i   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 95)) || ((sprite_column + 26 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�   �   �           �   h   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�i     �   g   i   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 95)) || ((sprite_column + 106 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�   �   �           �   m   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�n     �   l   n   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 13)) || ((sprite_column + 28 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�   �              �   m   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�r     �   l   n   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 13)) || ((sprite_column + 28 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�   �                m   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�z     �   l   n   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 13)) || ((sprite_column + 108 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�                  m   `    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�     �   l   n   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 93)) || ((sprite_column + 108 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�                 r   `    ����                                                                                                                                                                                                                                                                                                                            W           5           v        dÉ     �   q   s   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 30 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�                 r   a    ����                                                                                                                                                                                                                                                                                                                            W           5           v        dÌ     �   q   s   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column +80 < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 30 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�                 r   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        dÒ     �   q   s   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 11)) || ((sprite_column + 30 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�                 r   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        dÔ     �   q   s   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 191)) || ((sprite_column + 30 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�                 r   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        dÙ     �   q   s   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 91)) || ((sprite_column + 30 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�                 r   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        dë     �   q   s   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 91)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�    	             w   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        dñ     �   v   x   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 33) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 9)) || ((sprite_column + 32 < pixel_column) && (pixel_column < sprite_column + 41))))5�_�    
          	   w   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d÷     �   v   x   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 33) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 9)) || ((sprite_column + 32 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�  	            
   w   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        dý     �   v   x   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 33) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 9)) || ((sprite_column + 112 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�  
               w   `    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d��     �   v   x   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 33) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 89)) || ((sprite_column + 112 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�                         ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             z    else if ((pixel_row == sprite_row  + 1) && (sprite_column + 82 < pixel_column) && (pixel_column < sprite_column + 99))5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     begin5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             "            barrier_pix = 4'b1111;5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     end   5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                 // Row 2 5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             z    else if ((sprite_row + 2 == pixel_row) && (sprite_column + 81 < pixel_column) && (pixel_column < sprite_column + 100))5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     begin5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             "            barrier_pix = 4'b1111;5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     end   5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                 // Rows 3 - 9 5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             �    else if ((sprite_row + 2 < pixel_row) && (pixel_row < sprite_row  + 10) && (sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 101))5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     begin5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             "            barrier_pix = 4'b1111;5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     end5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                 // Row 105�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             �    else if ((sprite_row + 10 == pixel_row) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 88)) || ((sprite_column + 93 < pixel_column) && (pixel_column < sprite_column + 101))))5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     begin5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             "            barrier_pix = 4'b1111;5�_�                        ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     end5�_�                         ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                 // Row 11 5�_�    !                     ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             �    else if ((sprite_row + 11 == pixel_row) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 87)) || ((sprite_column + 94 < pixel_column) && (pixel_column < sprite_column + 101))))5�_�     "          !          ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     begin5�_�  !  #          "          ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             "            barrier_pix = 4'b1111;5�_�  "  $          #          ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     end5�_�  #  %          $          ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                 // Rows 12 & 135�_�  $  &          %          ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             �    else if ((sprite_row + 11 < pixel_row) && (pixel_row < sprite_row + 14) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 86)) || ((sprite_column + 95 < pixel_column) && (pixel_column < sprite_column + 101))))5�_�  %  '          &          ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     begin5�_�  &  (          '          ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             "            barrier_pix = 4'b1111;5�_�  '  )          (          ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     end5�_�  (  *          )          ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                 // Row 14, 15 and 16 5�_�  )  +          *          ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             �    else if ((sprite_row + 13 < pixel_row) && (pixel_row < sprite_row + 17) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 85)) || ((sprite_column + 96 < pixel_column) && (pixel_column < sprite_column + 101))))5�_�  *  ,          +          ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     begin5�_�  +  -          ,          ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~             "            barrier_pix = 4'b1111;5�_�  ,  .          -          ����                                                                                                                                                                                                                                                                                                                            {           W           v���    d��     �   ~                     end5�_�  -  /          .           ����                                                                                                                                                                                                                                                                                                                            {           Y           v        d��     �   ~   �   �       �      �   �    5�_�  .  0          /   |        ����                                                                                                                                                                                                                                                                                                                            {           Y           v        d��     �   {   |           5�_�  /  1          0   }       ����                                                                                                                                                                                                                                                                                                                            {           Y           v        d�     �   |   ~   �      9    // Row one of Barrier3's Sprite (Offset = 120 pix)   5�_�  0  2          1   }       ����                                                                                                                                                                                                                                                                                                                            {           Y           v        d�     �   |   ~   �      8    // Row ne of Barrier3's Sprite (Offset = 120 pix)   5�_�  1  3          2   }       ����                                                                                                                                                                                                                                                                                                                            {           Y           v        d�     �   |   ~   �      7    // Row e of Barrier3's Sprite (Offset = 120 pix)   5�_�  2  4          3   }       ����                                                                                                                                                                                                                                                                                                                            {           Y           v        d�
     �   |   ~   �      6    // Row  of Barrier3's Sprite (Offset = 120 pix)   5�_�  3  5          4   V       ����                                                                                                                                                                                                                                                                                                                            {           Y           v        d�     �   U   X   �              end5�_�  4  6          5   ~   2    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        d�%     �   }      �      ;    // Row 1 & 2 of Barrier3's Sprite (Offset = 120 pix)   5�_�  5  7          6      [    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        d�1     �   ~   �   �      �    else if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) && (sprite_column + 84 < pixel_column) && (pixel_column < sprite_column + 117))5�_�  6  8          7      �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        d�<     �   ~   �   �      �    else if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) && (sprite_column + 164 < pixel_column) && (pixel_column < sprite_column + 117))5�_�  7  9          8   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        d�L     �   �   �   �      �    else if ((sprite_row + 2 < pixel_row) && (pixel_row < sprite_row + 5) && (sprite_column + 82 < pixel_column) && (pixel_column < sprite_column + 119))5�_�  8  :          9   �   _    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        d�P     �   �   �   �      �    else if ((sprite_row + 2 < pixel_row) && (pixel_row < sprite_row + 5) && (sprite_column + 82 < pixel_column) && (pixel_column < sprite_column + 199))5�_�  9  ;          :   �   a    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        d�T     �   �   �   �      �    else if ((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) && (sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 121))5�_�  :  <          ;   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        d�X     �   �   �   �      �    else if ((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) && (sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 121))5�_�  ;  =          <   �   c    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        d�c     �   �   �   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 95)) || ((sprite_column + 106 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�  <  >          =   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        d�r     �   �   �   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 95)) || ((sprite_column + 106 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�  =  ?          >   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        d�w     �   �   �   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 175)) || ((sprite_column + 106 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�  >  @          ?   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        d�{     �   �   �   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 175)) || ((sprite_column + 186 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�  ?  A          @   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dĀ     �   �   �   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 93)) || ((sprite_column + 108 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�  @  B          A   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dĄ     �   �   �   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 93)) || ((sprite_column + 108 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  A  C          B   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dĊ     �   �   �   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 93)) || ((sprite_column + 188 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  B  D          C   �   c    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dď     �   �   �   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 173)) || ((sprite_column + 188 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  C  E          D   �   c    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dĒ     �   �   �   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 91)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�  D  F          E   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dĘ     �   �   �   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 91)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�  E  G          F   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dĞ     �   �   �   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 171)) || ((sprite_column + 110 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�  F  H          G   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dĢ     �   �   �   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 171)) || ((sprite_column + 190 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�  G  I          H   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dģ     �   �   �   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 171)) || ((sprite_column + 190 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�  H  J          I   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dħ     �   �   �   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 33) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 89)) || ((sprite_column + 112 < pixel_column) && (pixel_column < sprite_column + 121))))5�_�  I  K          J   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dĨ     �   �   �   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 33) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 89)) || ((sprite_column + 112 < pixel_column) && (pixel_column < sprite_column + 21))))5�_�  J  L          K   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dī     �   �   �   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 33) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 89)) || ((sprite_column + 112 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  K  M          L   �   �    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dı     �   �   �   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 33) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 89)) || ((sprite_column + 192 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  L  N          M   �   c    ����                                                                                                                                                                                                                                                                                                                            |           Z           v        dĸ     �   �   �   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 33) && (((sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 169)) || ((sprite_column + 192 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  M  O          N   �        ����                                                                                                                                                                                                                                                                                                                            �           �          v   !    d��     �   �   �   �   '               9    // Row one of Barrier4's Sprite (Offset = 120 pix)      |    else if ((pixel_row == sprite_row  + 1) && (sprite_column + 122 < pixel_column) && (pixel_column < sprite_column + 139))           begin   "            barrier_pix = 4'b1111;           end          // Row 2    {    else if ((sprite_row + 2 == pixel_row) && (sprite_column + 121 < pixel_column) && (pixel_column < sprite_column + 140))           begin   "            barrier_pix = 4'b1111;           end          // Rows 3 - 9    �    else if ((sprite_row + 2 < pixel_row) && (pixel_row < sprite_row  + 10) && (sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 141))           begin   "            barrier_pix = 4'b1111;           end       // Row 10   �    else if ((sprite_row + 10 == pixel_row) && (((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 128)) || ((sprite_column + 133 < pixel_column) && (pixel_column < sprite_column + 141))))           begin   "            barrier_pix = 4'b1111;           end       // Row 11    �    else if ((sprite_row + 11 == pixel_row) && (((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 127)) || ((sprite_column + 134 < pixel_column) && (pixel_column < sprite_column + 141))))           begin   "            barrier_pix = 4'b1111;           end       // Rows 12 & 13   �    else if ((sprite_row + 11 < pixel_row) && (pixel_row < sprite_row + 14) && (((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 126)) || ((sprite_column + 135 < pixel_column) && (pixel_column < sprite_column + 141))))           begin   "            barrier_pix = 4'b1111;           end       // Row 14, 15 and 16    �    else if ((sprite_row + 13 < pixel_row) && (pixel_row < sprite_row + 17) && (((sprite_column + 120 < pixel_column) && (pixel_column < sprite_column + 125)) || ((sprite_column + 136 < pixel_column) && (pixel_column < sprite_column + 141))))           begin   "            barrier_pix = 4'b1111;           end       else5�_�  N  P          O   �        ����                                                                                                                                                                                                                                                                                                                            �           �          v   !    d��     �   �   �   �          else5�_�  O  Q          P   �       ����                                                                                                                                                                                                                                                                                                                            �           �          v   !    d��     �   �   �   �              else5�_�  P  R          Q   �       ����                                                                                                                                                                                                                                                                                                                            �           �          v   !    d��     �   �   �   �       else5�_�  Q  S          R   �        ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d��     �   �   �   �          �   �   �   �    5�_�  R  T          S   �       ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d��     �   �   �   �      <     // Row 1 & 2 of Barrier3's Sprite (Offset = 160 pix)   5�_�  S  U          T   �       ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d��     �   �   �   �      ;    // Row 1 & 2 of Barrier3's Sprite (Offset = 160 pix)   5�_�  T  V          U   �   0    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d��     �   �   �   �      ;    // Row 1 & 2 of Barrier5's Sprite (Offset = 160 pix)   5�_�  U  W          V   �   0    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d��     �   �   �   �      :    // Row 1 & 2 of Barrier5's Sprite (Offset = 60 pix)   5�_�  V  X          W   �   0    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d��     �   �   �   �      9    // Row 1 & 2 of Barrier5's Sprite (Offset = 0 pix)   5�_�  W  Y          X   �   0    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d��     �   �   �   �      8    // Row 1 & 2 of Barrier5's Sprite (Offset =  pix)   5�_�  X  Z          Y   �   \    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d��     �   �   �   �      �    else if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) && (sprite_column + 164 < pixel_column) && (pixel_column < sprite_column + 197))5�_�  Y  [          Z   �   ^    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�      �   �   �   �      �    else if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) && (sprite_column + 2444 < pixel_column) && (pixel_column < sprite_column + 197))5�_�  Z  \          [   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�     �   �   �   �      �    else if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) && (sprite_column + 244 < pixel_column) && (pixel_column < sprite_column + 197))5�_�  [  ]          \   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�     �   �   �   �      �    else if ((sprite_row + 2 < pixel_row) && (pixel_row < sprite_row + 5) && (sprite_column + 162 < pixel_column) && (pixel_column < sprite_column + 199))5�_�  \  ^          ]   �   `    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�     �   �   �   �      �    else if ((sprite_row + 2 < pixel_row) && (pixel_row < sprite_row + 5) && (sprite_column + 162 < pixel_column) && (pixel_column < sprite_column + 279))5�_�  ]  _          ^   �   b    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�     �   �   �   �      �    else if ((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) && (sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 201))5�_�  ^  `          _   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�%     �   �   �   �      �    else if ((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) && (sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 201))5�_�  _  a          `   �   d    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�,     �   �   �   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 175)) || ((sprite_column + 186 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  `  b          a   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�9     �   �   �   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 175)) || ((sprite_column + 186 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  a  c          b   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�D     �   �   �   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 255)) || ((sprite_column + 186 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  b  d          c   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�I     �   �   �   �      �    else if ((sprite_row + 18 < pixel_row) && (pixel_row < sprite_row + 21) && (((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 255)) || ((sprite_column + 266 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  c  e          d   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�L     �   �   �   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 173)) || ((sprite_column + 188 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  d  f          e   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�P     �   �   �   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 173)) || ((sprite_column + 188 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  e  g          f   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�U     �   �   �   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 173)) || ((sprite_column + 268 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  f  h          g   �   d    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�Z     �   �   �   �      �    else if ((sprite_row + 20 < pixel_row) && (pixel_row < sprite_row + 23) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 253)) || ((sprite_column + 268 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  g  i          h   �   d    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�^     �   �   �   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 171)) || ((sprite_column + 190 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  h  j          i   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�c     �   �   �   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 171)) || ((sprite_column + 190 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  i  k          j   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�i     �   �   �   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 190 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  j  l          k   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�p     �   �   �   �      �    else if ((sprite_row + 22 < pixel_row) && (pixel_row < sprite_row + 27) && (((sprite_column + 240 < pixel_column) && (pixel_column < sprite_column + 251)) || ((sprite_column + 270 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  k  m          l   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�s     �   �   �   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 33) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 169)) || ((sprite_column + 192 < pixel_column) && (pixel_column < sprite_column + 201))))5�_�  l  n          m   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        d�y     �   �   �   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 33) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 169)) || ((sprite_column + 192 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  m  o          n   �   �    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        dń     �   �   �   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 33) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 169)) || ((sprite_column + 272 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  n  p          o   �   e    ����                                                                                                                                                                                                                                                                                                                            �           ~           v        dň     �   �   �   �      �    else if ((sprite_row + 26 < pixel_row) && (pixel_row < sprite_row + 33) && (((sprite_column + 160 < pixel_column) && (pixel_column < sprite_column + 249)) || ((sprite_column + 272 < pixel_column) && (pixel_column < sprite_column + 281))))5�_�  o  q          p   �        ����                                                                                                                                                                                                                                                                                                                            �           ~           v        dŎ     �   �   �   �              end    �   �   �   �       5�_�  p  r          q   �       ����                                                                                                                                                                                                                                                                                                                            �           ~           v        dŏ     �   �   �   �              end    �   �   �   �             �   �   �   �          5�_�  q  s          r   �       ����                                                                                                                                                                                                                                                                                                                            �           ~           v        dř     �   �   �   �      ;    // Row 1 & 2 of Barrier5's Sprite (Offset = 240 pix)   5�_�  r  t          s   �       ����                                                                                                                                                                                                                                                                                                                            �           ~           v        dŚ    �   �   �   �      <    // Row 1 & 2 of Barrierx5's Sprite (Offset = 240 pix)   5�_�  s  u          t   !       ����                                                                                                                                                                                                                                                                                                                                                             dɄ    �       "   �      <    // Initializing barriers 30 rows above the player sprite5�_�  t  v          u   #       ����                                                                                                                                                                                                                                                                                                                                                             dɩ     �   "   $   �          sprite_column = 250;5�_�  u  w          v   #       ����                                                                                                                                                                                                                                                                                                                                                             dɬ    �   "   $   �          sprite_column = 290;5�_�  v  x          w   !       ����                                                                                                                                                                                                                                                                                                                                                             d��     �       "   �      <    // Initializing barriers 40 rows above the player sprite5�_�  w  y          x   #       ����                                                                                                                                                                                                                                                                                                                                                             d��     �   "   $   �          sprite_column = 291;5�_�  x  z          y   #       ����                                                                                                                                                                                                                                                                                                                                                             d��     �   "   $   �          sprite_column = 91;5�_�  y  {          z   #       ����                                                                                                                                                                                                                                                                                                                                                             d��     �   "   $   �          sprite_column = 1;5�_�  z  |          {   #       ����                                                                                                                                                                                                                                                                                                                                                             d��     �   "   $   �          sprite_column = ;5�_�  {  }          |   $       ����                                                                                                                                                                                                                                                                                                                                                             d��     �   #   %   �          sprite_row = 430;5�_�  |  ~          }   "   5    ����                                                                                                                                                                                                                                                                                                                                                             d��     �   !   #   �      >    // and close to centered as possible. Columns: 251 <-> 3905�_�  }            ~   "   =    ����                                                                                                                                                                                                                                                                                                                                                             d�     �   !   #   �      >    // and close to centered as possible. Columns: 181 <-> 3905�_�  ~                 #       ����                                                                                                                                                                                                                                                                                                                                                             d�    �   "   $   �          sprite_column = 400;5�_�   �           �   �   c   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�B     �   b   d   �      �    else if ((sprite_row + 4 < pixel_row) && (pixel_row < sprite_row  + 19) && (sprite_column + 80 < pixel_column) && (pixel_column < sprite_column + 8u1))5�_�   �       �   �   �   Y   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�     �   X   Z   �      �    else if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) && (sprite_column + 84 < pixel_column) && (pixel_column < sprite_column + 7))5�_�   �           �   �   Y   �    ����                                                                                                                                                                                                                                                                                                                            W           5           v        d�     �   X   Z   �      �    else if ((sprite_row < pixel_row) && (pixel_row < sprite_row + 3) && (sprite_column + 84 < pixel_column) && (pixel_column < sprite_column + ))5�_�   �           �   �   Z        ����                                                                                                                                                                                                                                                                                                                            W           4           v        d��     �   Z   [   �    �   Z   [   �              end5�_�   a           c   b   D       ����                                                                                                                                                                                                                                                                                                                            5          5   @       v   @    d��     �   D   E   �    �   C   E   �      �    else if (((sprite_row + 10 == pixel_row) && (((sprite_column < pixel_column) && (pixel_column < sprite_column + 8)) || ((sprite_column + 13 < pixel_column) && (pixel_column < sprite_column + 21))))5��